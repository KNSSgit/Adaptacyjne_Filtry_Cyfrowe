//////////////////////////////////////////////////////////////////////////////////
// Kolo Naukowe Systemow Scalonych
// 10.2017
// 
// Modul: generator
// Projekt: Adaptacyjne filtry cyfrowe do kondycjonowania sygnalow biomedycznych 
// Model urzadzenia: Nexys Video Artix 7 (XC7A200T-1SBG484C)
// 
// Wersja: 0.1
//////////////////////////////////////////////////////////////////////////////////


module generator(
    output reg signed [23:0] data_out,
    input clk,
    input reset
    );
    
    reg signed [23:0] rom [0:399];
    reg [8:0] i;
    reg [15:0] counter;//5000 * 400pr�bek = 2 000 000 ; zegar 100mhz => 50hz

    always @(reset)
        begin
rom[0] = 24'b000000000000000000000000;
        rom[1] = 24'b000001000000011001011110;
        rom[2] = 24'b000010000000100111110001;
        rom[3] = 24'b000011000000011111110000;
        rom[4] = 24'b000011111111110110010111;
        rom[5] = 24'b000100111110100000101011;
        rom[6] = 24'b000101111100010011111011;
        rom[7] = 24'b000110111001000101100110;
        rom[8] = 24'b000111110100101011011000;
        rom[9] = 24'b001000101110111011010010;
        rom[10] = 24'b001001100111101011101000;
        rom[11] = 24'b001010011110110011000110;
        rom[12] = 24'b001011010100001000110011;
        rom[13] = 24'b001100000111100100010001;
        rom[14] = 24'b001100111000111101011111;
        rom[15] = 24'b001101101000001100111110;
        rom[16] = 24'b001110010101001011101110;
        rom[17] = 24'b001110111111110011010100;
        rom[18] = 24'b001111100111111101111010;
        rom[19] = 24'b010000001101100110010000;
        rom[20] = 24'b010000110000100111101101;
        rom[21] = 24'b010001010000111110010010;
        rom[22] = 24'b010001101110100110101001;
        rom[23] = 24'b010010001001011110000100;
        rom[24] = 24'b010010100001100010100100;
        rom[25] = 24'b010010110110110010110011;
        rom[26] = 24'b010011001001001110000111;
        rom[27] = 24'b010011011000110100100010;
        rom[28] = 24'b010011100101100110110000;
        rom[29] = 24'b010011101111100110001100;
        rom[30] = 24'b010011110110110100111001;
        rom[31] = 24'b010011111011010101100101;
        rom[32] = 24'b010011111101001011101000;
        rom[33] = 24'b010011111100011011000011;
        rom[34] = 24'b010011111001001000011110;
        rom[35] = 24'b010011110011011001001000;
        rom[36] = 24'b010011101011010010110011;
        rom[37] = 24'b010011100000111011111000;
        rom[38] = 24'b010011010100011011001111;
        rom[39] = 24'b010011000101111000010001;
        rom[40] = 24'b010010110101011010110100;
        rom[41] = 24'b010010100011001011001100;
        rom[42] = 24'b010010001111010010000110;
        rom[43] = 24'b010001111001111000100101;
        rom[44] = 24'b010001100011001000000011;
        rom[45] = 24'b010001001011001010001101;
        rom[46] = 24'b010000110010001000111110;
        rom[47] = 24'b010000011000001110100010;
        rom[48] = 24'b001111111101100101001101;
        rom[49] = 24'b001111100010010111011101;
        rom[50] = 24'b001111000110101111110110;
        rom[51] = 24'b001110101010111000111110;
        rom[52] = 24'b001110001110111101011011;
        rom[53] = 24'b001101110011000111110010;
        rom[54] = 24'b001101010111100010100010;
        rom[55] = 24'b001100111100011000000010;
        rom[56] = 24'b001100100001110010011101;
        rom[57] = 24'b001100000111111011110100;
        rom[58] = 24'b001011101110111101110110;
        rom[59] = 24'b001011010111000001111111;
        rom[60] = 24'b001011000000010001011000;
        rom[61] = 24'b001010101010110100110011;
        rom[62] = 24'b001010010110110100100111;
        rom[63] = 24'b001010000100011000110001;
        rom[64] = 24'b001001110011101000101111;
        rom[65] = 24'b001001100100101011100001;
        rom[66] = 24'b001001010111100111100101;
        rom[67] = 24'b001001001100100010110110;
        rom[68] = 24'b001001000011100010101010;
        rom[69] = 24'b001000111100101011110001;
        rom[70] = 24'b001000111000000010010110;
        rom[71] = 24'b001000110101101001111010;
        rom[72] = 24'b001000110101100101010011;
        rom[73] = 24'b001000110111110110110001;
        rom[74] = 24'b001000111100011111110111;
        rom[75] = 24'b001001000011100001011101;
        rom[76] = 24'b001001001100111011110001;
        rom[77] = 24'b001001011000101110010101;
        rom[78] = 24'b001001100110111000000000;
        rom[79] = 24'b001001110111010110111101;
        rom[80] = 24'b001010001010001000101110;
        rom[81] = 24'b001010011111001010001011;
        rom[82] = 24'b001010110110010111100001;
        rom[83] = 24'b001011001111101100010111;
        rom[84] = 24'b001011101011000011101100;
        rom[85] = 24'b001100001000010111111000;
        rom[86] = 24'b001100100111100010110001;
        rom[87] = 24'b001101001000011101101000;
        rom[88] = 24'b001101101011000001001101;
        rom[89] = 24'b001110001111000101110001;
        rom[90] = 24'b001110110100100011001000;
        rom[91] = 24'b001111011011010000101001;
        rom[92] = 24'b010000000011000101010100;
        rom[93] = 24'b010000101011110111101111;
        rom[94] = 24'b010001010101011110001110;
        rom[95] = 24'b010001111111101110110001;
        rom[96] = 24'b010010101010011111001010;
        rom[97] = 24'b010011010101100100111100;
        rom[98] = 24'b010100000000110101100000;
        rom[99] = 24'b010100101100000110001000;
        rom[100] = 24'b010101010111001100000000;
        rom[101] = 24'b010110000001111100010011;
        rom[102] = 24'b010110101100001100001010;
        rom[103] = 24'b010111010101110000110011;
        rom[104] = 24'b010111111110011111100001;
        rom[105] = 24'b011000100110001101110001;
        rom[106] = 24'b011001001100110001001000;
        rom[107] = 24'b011001110001111111011011;
        rom[108] = 24'b011010010101101110110001;
        rom[109] = 24'b011010110111110101100000;
        rom[110] = 24'b011011011000001010010101;
        rom[111] = 24'b011011110110100100010111;
        rom[112] = 24'b011100010010111011000101;
        rom[113] = 24'b011100101101000110011000;
        rom[114] = 24'b011101000100111110101011;
        rom[115] = 24'b011101011010011100110111;
        rom[116] = 24'b011101101101011010011000;
        rom[117] = 24'b011101111101110001001100;
        rom[118] = 24'b011110001011011011111000;
        rom[119] = 24'b011110010110010101100111;
        rom[120] = 24'b011110011110011010001011;
        rom[121] = 24'b011110100011100101111111;
        rom[122] = 24'b011110100101110110001001;
        rom[123] = 24'b011110100101001000011000;
        rom[124] = 24'b011110100001011011000111;
        rom[125] = 24'b011110011010101101011101;
        rom[126] = 24'b011110010000111111001101;
        rom[127] = 24'b011110000100010000110100;
        rom[128] = 24'b011101110100100011011100;
        rom[129] = 24'b011101100001111000111011;
        rom[130] = 24'b011101001100010011110011;
        rom[131] = 24'b011100110011110111001110;
        rom[132] = 24'b011100011000100111000001;
        rom[133] = 24'b011011111010100111101011;
        rom[134] = 24'b011011011001111110010010;
        rom[135] = 24'b011010110110110000100001;
        rom[136] = 24'b011010010001000100101001;
        rom[137] = 24'b011001101001000001100001;
        rom[138] = 24'b011000111110101110011111;
        rom[139] = 24'b011000010010010011011010;
        rom[140] = 24'b010111100011111000100110;
        rom[141] = 24'b010110110011100110110101;
        rom[142] = 24'b010110000001100111010010;
        rom[143] = 24'b010101001110000011100000;
        rom[144] = 24'b010100011001000101010111;
        rom[145] = 24'b010011100010110111000001;
        rom[146] = 24'b010010101011100010111010;
        rom[147] = 24'b010001110011010011101010;
        rom[148] = 24'b010000111010010100000101;
        rom[149] = 24'b010000000000101111001001;
        rom[150] = 24'b001111000110101111110110;
        rom[151] = 24'b001110001100100001010010;
        rom[152] = 24'b001101010010001110100011;
        rom[153] = 24'b001100011000000010101010;
        rom[154] = 24'b001011011110001000100111;
        rom[155] = 24'b001010100100101011001101;
        rom[156] = 24'b001001101011110101001010;
        rom[157] = 24'b001000110011110000111001;
        rom[158] = 24'b000111111100101000101001;
        rom[159] = 24'b000111000110100110010110;
        rom[160] = 24'b000110010001110011100111;
        rom[161] = 24'b000101011110011001101010;
        rom[162] = 24'b000100101100100001010111;
        rom[163] = 24'b000011111100010011001000;
        rom[164] = 24'b000011001101110110111001;
        rom[165] = 24'b000010100001010100001000;
        rom[166] = 24'b000001110110110001110010;
        rom[167] = 24'b000001001110010110001110;
        rom[168] = 24'b000000101000000111010001;
        rom[169] = 24'b000000000100001010001001;
        rom[170] = 24'b111111100010100011011101;
        rom[171] = 24'b111111000011010111001011;
        rom[172] = 24'b111110100110101000101000;
        rom[173] = 24'b111110001100011010011111;
        rom[174] = 24'b111101110100101110110001;
        rom[175] = 24'b111101011111100110110011;
        rom[176] = 24'b111101001101000011001111;
        rom[177] = 24'b111100111101000100000010;
        rom[178] = 24'b111100101111101000100000;
        rom[179] = 24'b111100100100101111010001;
        rom[180] = 24'b111100011100010110010001;
        rom[181] = 24'b111100010110011010110100;
        rom[182] = 24'b111100010010111001100010;
        rom[183] = 24'b111100010001101110011110;
        rom[184] = 24'b111100010010110101000001;
        rom[185] = 24'b111100010110000111111110;
        rom[186] = 24'b111100011011100001100101;
        rom[187] = 24'b111100100010111011100001;
        rom[188] = 24'b111100101100001110111011;
        rom[189] = 24'b111100110111010100100000;
        rom[190] = 24'b111101000100000100011010;
        rom[191] = 24'b111101010010010110011100;
        rom[192] = 24'b111101100010000001111100;
        rom[193] = 24'b111101110010111101111010;
        rom[194] = 24'b111110000101000001000010;
        rom[195] = 24'b111110011000000001101011;
        rom[196] = 24'b111110101011110101111111;
        rom[197] = 24'b111111000000010011111000;
        rom[198] = 24'b111111010101010001000111;
        rom[199] = 24'b111111101010100011010100;
        rom[200] = 24'b000000000000000000000000;
        rom[201] = 24'b000000010101011100101100;
        rom[202] = 24'b000000101010101110111001;
        rom[203] = 24'b000000111111101100001000;
        rom[204] = 24'b000001010100001010000001;
        rom[205] = 24'b000001100111111110010101;
        rom[206] = 24'b000001111010111110111110;
        rom[207] = 24'b000010001101000010000110;
        rom[208] = 24'b000010011101111110000100;
        rom[209] = 24'b000010101101101001100100;
        rom[210] = 24'b000010111011111011100110;
        rom[211] = 24'b000011001000101011100000;
        rom[212] = 24'b000011010011110001000101;
        rom[213] = 24'b000011011101000100011111;
        rom[214] = 24'b000011100100011110011011;
        rom[215] = 24'b000011101001111000000010;
        rom[216] = 24'b000011101101001010111111;
        rom[217] = 24'b000011101110010001100010;
        rom[218] = 24'b000011101101000110011110;
        rom[219] = 24'b000011101001100101001100;
        rom[220] = 24'b000011100011101001101111;
        rom[221] = 24'b000011011011010000101111;
        rom[222] = 24'b000011010000010111100000;
        rom[223] = 24'b000011000010111011111110;
        rom[224] = 24'b000010110010111100110001;
        rom[225] = 24'b000010100000011001001101;
        rom[226] = 24'b000010001011010001001111;
        rom[227] = 24'b000001110011100101100001;
        rom[228] = 24'b000001011001010111011000;
        rom[229] = 24'b000000111100101000110101;
        rom[230] = 24'b000000011101011100100011;
        rom[231] = 24'b111111111011110101110111;
        rom[232] = 24'b111111010111111000101111;
        rom[233] = 24'b111110110001101001110010;
        rom[234] = 24'b111110001001001110001110;
        rom[235] = 24'b111101011110101011111000;
        rom[236] = 24'b111100110010001001000111;
        rom[237] = 24'b111100000011101100111000;
        rom[238] = 24'b111011010011011110101001;
        rom[239] = 24'b111010100001100110010110;
        rom[240] = 24'b111001101110001100011001;
        rom[241] = 24'b111000111001011001101010;
        rom[242] = 24'b111000000011010111010111;
        rom[243] = 24'b110111001100001111000111;
        rom[244] = 24'b110110010100001010110110;
        rom[245] = 24'b110101011011010100110011;
        rom[246] = 24'b110100100001110111011001;
        rom[247] = 24'b110011100111111101010110;
        rom[248] = 24'b110010101101110001011101;
        rom[249] = 24'b110001110011011110101110;
        rom[250] = 24'b110000111001010000001010;
        rom[251] = 24'b101111111111010000110111;
        rom[252] = 24'b101111000101101011111011;
        rom[253] = 24'b101110001100101100010110;
        rom[254] = 24'b101101010100011101000110;
        rom[255] = 24'b101100011101001000111111;
        rom[256] = 24'b101011100110111010101001;
        rom[257] = 24'b101010110001111100100000;
        rom[258] = 24'b101001111110011000101110;
        rom[259] = 24'b101001001100011001001011;
        rom[260] = 24'b101000011100000111011010;
        rom[261] = 24'b100111101101101100100110;
        rom[262] = 24'b100111000001010001100001;
        rom[263] = 24'b100110010110111110011111;
        rom[264] = 24'b100101101110111011010111;
        rom[265] = 24'b100101001001001111011111;
        rom[266] = 24'b100100100110000001101110;
        rom[267] = 24'b100100000101011000010101;
        rom[268] = 24'b100011100111011000111111;
        rom[269] = 24'b100011001100001000110010;
        rom[270] = 24'b100010110011101100001101;
        rom[271] = 24'b100010011110000111000101;
        rom[272] = 24'b100010001011011100100100;
        rom[273] = 24'b100001111011101111001100;
        rom[274] = 24'b100001101111000000110011;
        rom[275] = 24'b100001100101010010100011;
        rom[276] = 24'b100001011110100100111001;
        rom[277] = 24'b100001011010110111101000;
        rom[278] = 24'b100001011010001001110111;
        rom[279] = 24'b100001011100011010000001;
        rom[280] = 24'b100001100001100101110101;
        rom[281] = 24'b100001101001101010011001;
        rom[282] = 24'b100001110100100100001000;
        rom[283] = 24'b100010000010001110110100;
        rom[284] = 24'b100010010010100101101000;
        rom[285] = 24'b100010100101100011001001;
        rom[286] = 24'b100010111011000001010101;
        rom[287] = 24'b100011010010111001101000;
        rom[288] = 24'b100011101101000100111011;
        rom[289] = 24'b100100001001011011101001;
        rom[290] = 24'b100100100111110101101011;
        rom[291] = 24'b100101001000001010100000;
        rom[292] = 24'b100101101010010001001111;
        rom[293] = 24'b100110001110000000100101;
        rom[294] = 24'b100110110011001110111000;
        rom[295] = 24'b100111011001110010001111;
        rom[296] = 24'b101000000001100000011111;
        rom[297] = 24'b101000101010001111001101;
        rom[298] = 24'b101001010011110011110110;
        rom[299] = 24'b101001111110000011101101;
        rom[300] = 24'b101010101000110100000000;
        rom[301] = 24'b101011010011111001111000;
        rom[302] = 24'b101011111111001010100000;
        rom[303] = 24'b101100101010011011000100;
        rom[304] = 24'b101101010101100000110110;
        rom[305] = 24'b101110000000010001001111;
        rom[306] = 24'b101110101010100001110010;
        rom[307] = 24'b101111010100001000010001;
        rom[308] = 24'b101111111100111010101100;
        rom[309] = 24'b110000100100101111010111;
        rom[310] = 24'b110001001011011100111000;
        rom[311] = 24'b110001110000111010001111;
        rom[312] = 24'b110010010100111110110011;
        rom[313] = 24'b110010110111100010011000;
        rom[314] = 24'b110011011000011101001111;
        rom[315] = 24'b110011110111101000001000;
        rom[316] = 24'b110100010100111100010100;
        rom[317] = 24'b110100110000010011101001;
        rom[318] = 24'b110101001001101000011111;
        rom[319] = 24'b110101100000110101110101;
        rom[320] = 24'b110101110101110111010010;
        rom[321] = 24'b110110001000101001000011;
        rom[322] = 24'b110110011001001000000000;
        rom[323] = 24'b110110100111010001101011;
        rom[324] = 24'b110110110011000100001111;
        rom[325] = 24'b110110111100011110100011;
        rom[326] = 24'b110111000011100000001001;
        rom[327] = 24'b110111001000001001001111;
        rom[328] = 24'b110111001010011010101101;
        rom[329] = 24'b110111001010010110000110;
        rom[330] = 24'b110111000111111101101010;
        rom[331] = 24'b110111000011010100001111;
        rom[332] = 24'b110110111100011101010110;
        rom[333] = 24'b110110110011011101001010;
        rom[334] = 24'b110110101000011000011011;
        rom[335] = 24'b110110011011010100011111;
        rom[336] = 24'b110110001100010111010001;
        rom[337] = 24'b110101111011100111001111;
        rom[338] = 24'b110101101001001011011001;
        rom[339] = 24'b110101010101001011001101;
        rom[340] = 24'b110100111111101110101000;
        rom[341] = 24'b110100101000111110000001;
        rom[342] = 24'b110100010001000010001010;
        rom[343] = 24'b110011111000000100001100;
        rom[344] = 24'b110011011110001101100011;
        rom[345] = 24'b110011000011100111111110;
        rom[346] = 24'b110010101000011101011110;
        rom[347] = 24'b110010001100111000001110;
        rom[348] = 24'b110001110001000010100101;
        rom[349] = 24'b110001010101000111000010;
        rom[350] = 24'b110000111001010000001010;
        rom[351] = 24'b110000011101101000100011;
        rom[352] = 24'b110000000010011010110011;
        rom[353] = 24'b101111100111110001011110;
        rom[354] = 24'b101111001101110111000010;
        rom[355] = 24'b101110110100110101110011;
        rom[356] = 24'b101110011100110111111101;
        rom[357] = 24'b101110000110000111011011;
        rom[358] = 24'b101101110000101101111010;
        rom[359] = 24'b101101011100110100110100;
        rom[360] = 24'b101101001010100101001100;
        rom[361] = 24'b101100111010000111101111;
        rom[362] = 24'b101100101011100100110001;
        rom[363] = 24'b101100011111000100001000;
        rom[364] = 24'b101100010100101101001101;
        rom[365] = 24'b101100001100100110111000;
        rom[366] = 24'b101100000110110111100010;
        rom[367] = 24'b101100000011100100111101;
        rom[368] = 24'b101100000010110100011000;
        rom[369] = 24'b101100000100101010011011;
        rom[370] = 24'b101100001001001011000111;
        rom[371] = 24'b101100010000011001110100;
        rom[372] = 24'b101100011010011001010000;
        rom[373] = 24'b101100100111001011011110;
        rom[374] = 24'b101100110110110001111001;
        rom[375] = 24'b101101001001001101001101;
        rom[376] = 24'b101101011110011101011100;
        rom[377] = 24'b101101110110100001111100;
        rom[378] = 24'b101110010001011001010111;
        rom[379] = 24'b101110101111000001101110;
        rom[380] = 24'b101111001111011000010011;
        rom[381] = 24'b101111110010011001110000;
        rom[382] = 24'b110000011000000010000110;
        rom[383] = 24'b110001000000001100101100;
        rom[384] = 24'b110001101010110100010010;
        rom[385] = 24'b110010010111110011000010;
        rom[386] = 24'b110011000111000010100001;
        rom[387] = 24'b110011111000011011101111;
        rom[388] = 24'b110100101011110111001101;
        rom[389] = 24'b110101100001001100111010;
        rom[390] = 24'b110110011000010100011000;
        rom[391] = 24'b110111010001000100101110;
        rom[392] = 24'b111000001011010100101000;
        rom[393] = 24'b111001000110111010011010;
        rom[394] = 24'b111010000011101100000101;
        rom[395] = 24'b111011000001011111010101;
        rom[396] = 24'b111100000000001001101001;
        rom[397] = 24'b111100111111100000010000;
        rom[398] = 24'b111101111111011000001111;
        rom[399] = 24'b111110111111100110100010;

        end
        
        always @(posedge(clk))
            begin
                if(reset)
                    begin
                        data_out <= 24'b0;
                        i <= 9'b0;
                        counter <= 16'b0;
                    end
                else
                    begin
                        if(counter == 16'd5000)
                            begin
                                data_out <= rom[i];
                                counter <= 16'b0;
                                if(i == 399) i <= 0;
                                else i <= i + 1;
                            end
                        else counter <= counter + 16'd1;
                    end
            end
            
endmodule
