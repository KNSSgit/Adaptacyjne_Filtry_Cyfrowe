module gen_ekg_60(
 	 output reg signed [23:0] data_out,
	 input clk,
	 input reset
	 ); 

	 reg signed [23:0] rom[0:1999];
	 reg [15:0] i;
	 reg [15:0] counter;//5000 * 2000pr�bek = 10 000 000 ; zegar 10mhz => 1hz

	 always @(reset)     // fs = 2kHz; f1 = 1Hz; A1 = 3000000; f2 = 60Hz; A2 = 90000
		 begin 
         rom[0] = 24'b111111110101110110001110;
         rom[1] = 24'b000000000100010100101101;
         rom[2] = 24'b000000001111010111010010;
         rom[3] = 24'b000000010000011100111100;
         rom[4] = 24'b000000011001111000000100;
         rom[5] = 24'b000000010010110001010000;
         rom[6] = 24'b000000010110010001000100;
         rom[7] = 24'b000000101000100100011010;
         rom[8] = 24'b000000011111010010001101;
         rom[9] = 24'b000000011010110100011101;
         rom[10] = 24'b000000101010011001000010;
         rom[11] = 24'b000000100111111111101101;
         rom[12] = 24'b000000011001001000101100;
         rom[13] = 24'b000000011000000111110110;
         rom[14] = 24'b000000100100100100011000;
         rom[15] = 24'b000000000101110001010010;
         rom[16] = 24'b000000000100000001101001;
         rom[17] = 24'b111111111110100001000011;
         rom[18] = 24'b111111110010110010110110;
         rom[19] = 24'b111111110011000011100000;
         rom[20] = 24'b111111100010100100000110;
         rom[21] = 24'b111111100000101111011011;
         rom[22] = 24'b111111100011010000110011;
         rom[23] = 24'b111111001100011001110101;
         rom[24] = 24'b111111011111110010100100;
         rom[25] = 24'b111111011001110001101101;
         rom[26] = 24'b111111010000001001100011;
         rom[27] = 24'b111111011000001101110101;
         rom[28] = 24'b111111010111111001101001;
         rom[29] = 24'b111111101001001010000100;
         rom[30] = 24'b111111101110100101000101;
         rom[31] = 24'b111111110110001001001000;
         rom[32] = 24'b111111110111011101110100;
         rom[33] = 24'b111111111111101111111001;
         rom[34] = 24'b000000001101100111000010;
         rom[35] = 24'b000000000011110110111111;
         rom[36] = 24'b000000011001111011101010;
         rom[37] = 24'b000000010100011101000011;
         rom[38] = 24'b000000100000101111100000;
         rom[39] = 24'b000000011001100010111110;
         rom[40] = 24'b000000011000111000111001;
         rom[41] = 24'b000000100111100110011011;
         rom[42] = 24'b000000100001011100000100;
         rom[43] = 24'b000000100000010000100100;
         rom[44] = 24'b000000100010001011100111;
         rom[45] = 24'b000000100100100111001110;
         rom[46] = 24'b000000001011000110110111;
         rom[47] = 24'b000000010001110010001110;
         rom[48] = 24'b111111111101001100100101;
         rom[49] = 24'b000000010111111011100011;
         rom[50] = 24'b111111111010110111110000;
         rom[51] = 24'b111111111000111011011100;
         rom[52] = 24'b111111111101001101100001;
         rom[53] = 24'b111111100100110010101011;
         rom[54] = 24'b111111110001101000101111;
         rom[55] = 24'b111111100011010110101010;
         rom[56] = 24'b111111011111011101001110;
         rom[57] = 24'b111111100000011000111001;
         rom[58] = 24'b111111010101110010111100;
         rom[59] = 24'b111111100111111100011101;
         rom[60] = 24'b111111010111011111011010;
         rom[61] = 24'b111111011100010000000001;
         rom[62] = 24'b111111101111100110110110;
         rom[63] = 24'b111111011101010010100011;
         rom[64] = 24'b111111101011110011010011;
         rom[65] = 24'b111111111010110111101101;
         rom[66] = 24'b111111101011011000011010;
         rom[67] = 24'b111111111100011010101101;
         rom[68] = 24'b000000001000111110111100;
         rom[69] = 24'b000000001110011111101101;
         rom[70] = 24'b000000001110110011010100;
         rom[71] = 24'b000000101000100010101000;
         rom[72] = 24'b000000011101000100000000;
         rom[73] = 24'b000000100011001001011001;
         rom[74] = 24'b000000100111000100001110;
         rom[75] = 24'b000000101011000001110101;
         rom[76] = 24'b000000101010111011001101;
         rom[77] = 24'b000000100011111010110101;
         rom[78] = 24'b000000100111010010101001;
         rom[79] = 24'b000000011110010000100011;
         rom[80] = 24'b000000010001111010111111;
         rom[81] = 24'b000000001101000000101001;
         rom[82] = 24'b000000000011000100101110;
         rom[83] = 24'b000000010001100010101001;
         rom[84] = 24'b111111111011001111000010;
         rom[85] = 24'b111111110010111111110011;
         rom[86] = 24'b111111101011001110101100;
         rom[87] = 24'b111111101011001011100011;
         rom[88] = 24'b111111100110011111000100;
         rom[89] = 24'b111111101111011111100000;
         rom[90] = 24'b111111011001010000100011;
         rom[91] = 24'b111111011000110100100110;
         rom[92] = 24'b111111100001001110001101;
         rom[93] = 24'b111111010110001010110001;
         rom[94] = 24'b111111100001101000101001;
         rom[95] = 24'b111111011110101001010000;
         rom[96] = 24'b111111101011101101111101;
         rom[97] = 24'b000000000001010010001101;
         rom[98] = 24'b111111101111000101011010;
         rom[99] = 24'b111111111010111001111111;
         rom[100] = 24'b000000000110000010100110;
         rom[101] = 24'b000000001001001111000001;
         rom[102] = 24'b000000000010000110100101;
         rom[103] = 24'b000000001000100111110000;
         rom[104] = 24'b000000011010110010111100;
         rom[105] = 24'b000000010110111011010000;
         rom[106] = 24'b000000011111011111101110;
         rom[107] = 24'b000000100010100101100100;
         rom[108] = 24'b000000110100110011110010;
         rom[109] = 24'b000000111001000100000010;
         rom[110] = 24'b000000011101011101010111;
         rom[111] = 24'b000000001111010011001010;
         rom[112] = 24'b000000100110001001011010;
         rom[113] = 24'b000000000101110101111110;
         rom[114] = 24'b000000001001111101101101;
         rom[115] = 24'b000000001101001111001001;
         rom[116] = 24'b111111110111101000100110;
         rom[117] = 24'b000000000111101110001010;
         rom[118] = 24'b111111101101001100000000;
         rom[119] = 24'b111111110001000111101000;
         rom[120] = 24'b111111101101010000010101;
         rom[121] = 24'b111111010001010111001010;
         rom[122] = 24'b111111010111000011101101;
         rom[123] = 24'b111111010011001001100110;
         rom[124] = 24'b111111011010000011001000;
         rom[125] = 24'b111111011000111110110111;
         rom[126] = 24'b111111010011011010011010;
         rom[127] = 24'b111111011011111011000111;
         rom[128] = 24'b111111010010101010011001;
         rom[129] = 24'b111111100001010100110110;
         rom[130] = 24'b111111101110000001010000;
         rom[131] = 24'b111111110111010110110011;
         rom[132] = 24'b111111110011101010011010;
         rom[133] = 24'b000000000111110001000111;
         rom[134] = 24'b000000000000011010100000;
         rom[135] = 24'b000000010000011011000101;
         rom[136] = 24'b000000010001111011100000;
         rom[137] = 24'b000000010100110111110011;
         rom[138] = 24'b000000100001000101100011;
         rom[139] = 24'b000000100000111010110011;
         rom[140] = 24'b000000101001101000101100;
         rom[141] = 24'b000000110001010110101110;
         rom[142] = 24'b000000010101100100011100;
         rom[143] = 24'b000000110000000001000110;
         rom[144] = 24'b000000100000110101010001;
         rom[145] = 24'b000000011110100011010110;
         rom[146] = 24'b000000010010111010111100;
         rom[147] = 24'b000000001111100110101001;
         rom[148] = 24'b000000010010000111011110;
         rom[149] = 24'b000000000010010000000111;
         rom[150] = 24'b111111111101110101111001;
         rom[151] = 24'b111111111001111010011111;
         rom[152] = 24'b111111100000100011100111;
         rom[153] = 24'b111111110100100100100110;
         rom[154] = 24'b111111101011011111001000;
         rom[155] = 24'b111111011001110000111100;
         rom[156] = 24'b111111001010000000010101;
         rom[157] = 24'b111111100001100010010000;
         rom[158] = 24'b111111010011011000001110;
         rom[159] = 24'b111111011000111010100001;
         rom[160] = 24'b111111011001111100001101;
         rom[161] = 24'b111111010000100011000101;
         rom[162] = 24'b111111100010011110010001;
         rom[163] = 24'b111111100110010010000111;
         rom[164] = 24'b111111110011000010000010;
         rom[165] = 24'b111111110001101000000001;
         rom[166] = 24'b111111111000000000111010;
         rom[167] = 24'b111111111111011111110100;
         rom[168] = 24'b000000000010110001000101;
         rom[169] = 24'b000000010001010100101100;
         rom[170] = 24'b000000010100011100011000;
         rom[171] = 24'b000000010101001001001110;
         rom[172] = 24'b000000101111010010010010;
         rom[173] = 24'b000000100011100011110011;
         rom[174] = 24'b000000100000100110100100;
         rom[175] = 24'b000000100110100010101000;
         rom[176] = 24'b000000101110111000000011;
         rom[177] = 24'b000000011000010110111011;
         rom[178] = 24'b000000001111110100001101;
         rom[179] = 24'b000000011111111010000111;
         rom[180] = 24'b000000010000010000001000;
         rom[181] = 24'b000000010111001011101100;
         rom[182] = 24'b111111111100010001001101;
         rom[183] = 24'b111111111101001101101001;
         rom[184] = 24'b000000000000101111101010;
         rom[185] = 24'b111111101111000110010100;
         rom[186] = 24'b111111101001011010100110;
         rom[187] = 24'b111111100101001101101110;
         rom[188] = 24'b111111101011001000100000;
         rom[189] = 24'b111111011011011010110110;
         rom[190] = 24'b111111010111001011100100;
         rom[191] = 24'b111111011000110111010010;
         rom[192] = 24'b111111011011011110001000;
         rom[193] = 24'b111111011010100001110110;
         rom[194] = 24'b111111100100100110111001;
         rom[195] = 24'b111111011111011100000001;
         rom[196] = 24'b111111100111000110011100;
         rom[197] = 24'b111111101000111001100010;
         rom[198] = 24'b111111111001111010000100;
         rom[199] = 24'b000000000000100101101000;
         rom[200] = 24'b000000001001100101101011;
         rom[201] = 24'b000000000010101101110000;
         rom[202] = 24'b000000001010011110111000;
         rom[203] = 24'b000000100011010101010111;
         rom[204] = 24'b000000010010111101110111;
         rom[205] = 24'b000000010010100110010010;
         rom[206] = 24'b000000011101011110010001;
         rom[207] = 24'b000000101001100010001010;
         rom[208] = 24'b000000011000101111101100;
         rom[209] = 24'b000000100101001001000001;
         rom[210] = 24'b000000011110000111101111;
         rom[211] = 24'b000000101001000111100011;
         rom[212] = 24'b000000010110110111010111;
         rom[213] = 24'b000000001011010001110101;
         rom[214] = 24'b000000011000011101111001;
         rom[215] = 24'b000000011010001010011000;
         rom[216] = 24'b000000000000110001010111;
         rom[217] = 24'b111111110111001110000000;
         rom[218] = 24'b000000000001100101010110;
         rom[219] = 24'b111111100101000111001000;
         rom[220] = 24'b111111110011010010001010;
         rom[221] = 24'b111111011100011110101110;
         rom[222] = 24'b111111110100010101110000;
         rom[223] = 24'b111111010001111101001101;
         rom[224] = 24'b111111011101011011010111;
         rom[225] = 24'b111111011001100101111111;
         rom[226] = 24'b111111011000010011000110;
         rom[227] = 24'b111111011011111000111001;
         rom[228] = 24'b111111101000010100110100;
         rom[229] = 24'b111111100001010001010010;
         rom[230] = 24'b111111110000010000111011;
         rom[231] = 24'b111111111010101000110100;
         rom[232] = 24'b111111110111100101111000;
         rom[233] = 24'b111111111111001011100101;
         rom[234] = 24'b111111111111010010000100;
         rom[235] = 24'b000000001101111010100100;
         rom[236] = 24'b000000001001011001010101;
         rom[237] = 24'b000000011111100010111011;
         rom[238] = 24'b000000010100010111100100;
         rom[239] = 24'b000000011001110101110100;
         rom[240] = 24'b000000101000011000010110;
         rom[241] = 24'b000000100011111001111010;
         rom[242] = 24'b000000100011000011010001;
         rom[243] = 24'b000000100101101011000011;
         rom[244] = 24'b000000100010000000111001;
         rom[245] = 24'b000000010100011001101000;
         rom[246] = 24'b000000100101010010001100;
         rom[247] = 24'b000000001000001100111010;
         rom[248] = 24'b000000010010010010001010;
         rom[249] = 24'b000000001011101100110101;
         rom[250] = 24'b111111111111001010110000;
         rom[251] = 24'b111111110110101010010100;
         rom[252] = 24'b111111101101100110111111;
         rom[253] = 24'b111111010110110110110010;
         rom[254] = 24'b111111110010110011000001;
         rom[255] = 24'b111111100110000100010000;
         rom[256] = 24'b111111100101011001010000;
         rom[257] = 24'b111111010101101011001010;
         rom[258] = 24'b111111101010110101111000;
         rom[259] = 24'b111111100101100010110011;
         rom[260] = 24'b111111100110110111011110;
         rom[261] = 24'b111111011111101010111111;
         rom[262] = 24'b111111100010100101000100;
         rom[263] = 24'b111111101110101010011110;
         rom[264] = 24'b111111101011010100000110;
         rom[265] = 24'b111111110100000101010110;
         rom[266] = 24'b111111110101100010100000;
         rom[267] = 24'b111111111011011000010101;
         rom[268] = 24'b000000000011010011111010;
         rom[269] = 24'b000000010001100010100000;
         rom[270] = 24'b000000011100111011101110;
         rom[271] = 24'b000000011111000110010100;
         rom[272] = 24'b000000100010110010111110;
         rom[273] = 24'b000000011000100001100101;
         rom[274] = 24'b000000101001000000010001;
         rom[275] = 24'b000000100110100100000100;
         rom[276] = 24'b000000101111011101110000;
         rom[277] = 24'b000000011110100101010001;
         rom[278] = 24'b000000110000100010010101;
         rom[279] = 24'b000000101001011001010101;
         rom[280] = 24'b000000010111110011111110;
         rom[281] = 24'b000000001100100100111111;
         rom[282] = 24'b000000010001011010010110;
         rom[283] = 24'b000000000101001010111010;
         rom[284] = 24'b111111110001010001000011;
         rom[285] = 24'b111111110100110110111110;
         rom[286] = 24'b111111111000100101101111;
         rom[287] = 24'b111111100011110001000000;
         rom[288] = 24'b111111101110000101100110;
         rom[289] = 24'b111111100100001001101000;
         rom[290] = 24'b111111101100110001011010;
         rom[291] = 24'b111111010111101001100000;
         rom[292] = 24'b111111100010011001000010;
         rom[293] = 24'b111111011101011101010111;
         rom[294] = 24'b111111001101101101111011;
         rom[295] = 24'b111111100011101011110011;
         rom[296] = 24'b111111101010011001000000;
         rom[297] = 24'b111111110000100000110110;
         rom[298] = 24'b111111110101000100011111;
         rom[299] = 24'b111111111001000011001001;
         rom[300] = 24'b000000000000000011100111;
         rom[301] = 24'b000000001000110011011010;
         rom[302] = 24'b000000001011010011011000;
         rom[303] = 24'b000000011000110001001111;
         rom[304] = 24'b000000010110001101010101;
         rom[305] = 24'b000000011110010010010011;
         rom[306] = 24'b000000100110110110000101;
         rom[307] = 24'b000000011100111000101110;
         rom[308] = 24'b000000100101011100001001;
         rom[309] = 24'b000000010001001001110101;
         rom[310] = 24'b000000011111100100111100;
         rom[311] = 24'b000000011011010111100111;
         rom[312] = 24'b000000011011110111001000;
         rom[313] = 24'b000000010010011001000111;
         rom[314] = 24'b000000001111001101001111;
         rom[315] = 24'b000000000111100011001011;
         rom[316] = 24'b000000000011101110011010;
         rom[317] = 24'b000000001100111011110010;
         rom[318] = 24'b111111110011110100110111;
         rom[319] = 24'b111111110111110000110010;
         rom[320] = 24'b111111100010010011101000;
         rom[321] = 24'b111111101110011011010111;
         rom[322] = 24'b111111010111111110000100;
         rom[323] = 24'b111111100100011011011101;
         rom[324] = 24'b111111010101101100101011;
         rom[325] = 24'b111111011000111011000011;
         rom[326] = 24'b111111011011011011000000;
         rom[327] = 24'b111111011110011111000100;
         rom[328] = 24'b111111010101011111000010;
         rom[329] = 24'b111111101001001010100111;
         rom[330] = 24'b111111110010100000001011;
         rom[331] = 24'b111111101011011100100100;
         rom[332] = 24'b111111110010000000111110;
         rom[333] = 24'b000000000010111000101000;
         rom[334] = 24'b000000000111100001011001;
         rom[335] = 24'b000000001001001010011100;
         rom[336] = 24'b000000010000011000110100;
         rom[337] = 24'b000000100101000101100001;
         rom[338] = 24'b000000010110001100100101;
         rom[339] = 24'b000000100001001101000101;
         rom[340] = 24'b000000100011110101010111;
         rom[341] = 24'b000000101000110011010001;
         rom[342] = 24'b000000101111100010001101;
         rom[343] = 24'b000000011110111010001100;
         rom[344] = 24'b000000011100011000101001;
         rom[345] = 24'b000000010100000101010111;
         rom[346] = 24'b000000001110100111001101;
         rom[347] = 24'b000000001010110110010000;
         rom[348] = 24'b000000001001000101110000;
         rom[349] = 24'b000000000101100101000110;
         rom[350] = 24'b000000000111010011100101;
         rom[351] = 24'b111111101101111001010111;
         rom[352] = 24'b111111110111111100111001;
         rom[353] = 24'b111111110010111001110000;
         rom[354] = 24'b111111100110001110011011;
         rom[355] = 24'b111111011110000011010101;
         rom[356] = 24'b111111100110100001100010;
         rom[357] = 24'b111111010110110001100100;
         rom[358] = 24'b111111100000010110101100;
         rom[359] = 24'b111111011001101111000010;
         rom[360] = 24'b111111011010111110101100;
         rom[361] = 24'b111111011100010010000001;
         rom[362] = 24'b111111011001101001101010;
         rom[363] = 24'b111111101001111010010000;
         rom[364] = 24'b111111110101011110100111;
         rom[365] = 24'b111111111010110000011011;
         rom[366] = 24'b111111111010101001100110;
         rom[367] = 24'b000000001010111010010110;
         rom[368] = 24'b111111110111010000111111;
         rom[369] = 24'b000000001100101111111111;
         rom[370] = 24'b000000010010100101010111;
         rom[371] = 24'b000000101010101111011111;
         rom[372] = 24'b000000100000100100011000;
         rom[373] = 24'b000000011000001001110010;
         rom[374] = 24'b000000100111110111101010;
         rom[375] = 24'b000000101000101001000110;
         rom[376] = 24'b000000011101110101110001;
         rom[377] = 24'b000000101010100001100110;
         rom[378] = 24'b000000100000000001101110;
         rom[379] = 24'b000000100000100110011010;
         rom[380] = 24'b000000010101011110010010;
         rom[381] = 24'b000000011011000011010111;
         rom[382] = 24'b000000001100101001011110;
         rom[383] = 24'b000000000001011111100100;
         rom[384] = 24'b111111111000101100111001;
         rom[385] = 24'b111111110111011100110011;
         rom[386] = 24'b111111110010000001101001;
         rom[387] = 24'b111111011110100001100110;
         rom[388] = 24'b111111101000010011010010;
         rom[389] = 24'b111111100000010001001001;
         rom[390] = 24'b111111100011010010111110;
         rom[391] = 24'b111111011011110011101010;
         rom[392] = 24'b111111100010010011001110;
         rom[393] = 24'b111111100010000110100110;
         rom[394] = 24'b111111100111101010010000;
         rom[395] = 24'b111111011111110000100100;
         rom[396] = 24'b111111110101110001010011;
         rom[397] = 24'b111111100100010010011110;
         rom[398] = 24'b111111111101011000110110;
         rom[399] = 24'b000000000010011000010010;
         rom[400] = 24'b000000000001000101110011;
         rom[401] = 24'b000000000001101011110111;
         rom[402] = 24'b000000010100000001001001;
         rom[403] = 24'b000000000010101010000011;
         rom[404] = 24'b000000100011001110101111;
         rom[405] = 24'b000000100001101110110111;
         rom[406] = 24'b000000010110111000010011;
         rom[407] = 24'b000000100111010001100010;
         rom[408] = 24'b000000101101101110010101;
         rom[409] = 24'b000000010010111101100111;
         rom[410] = 24'b000000100101101110000101;
         rom[411] = 24'b000000011011111001111100;
         rom[412] = 24'b000000011110100001001000;
         rom[413] = 24'b000000011011000000010111;
         rom[414] = 24'b000000001100111010001101;
         rom[415] = 24'b000000001000101111110101;
         rom[416] = 24'b000000000001101101110001;
         rom[417] = 24'b111111110101011100111111;
         rom[418] = 24'b000000000000000011111110;
         rom[419] = 24'b111111011101100000111010;
         rom[420] = 24'b111111100010011111001010;
         rom[421] = 24'b111111100010000001000101;
         rom[422] = 24'b111111101010000100101001;
         rom[423] = 24'b111111011100111011100110;
         rom[424] = 24'b111111011100100100000111;
         rom[425] = 24'b111111011100100011101110;
         rom[426] = 24'b111111010101110011000010;
         rom[427] = 24'b111111011111110110000011;
         rom[428] = 24'b111111100111011101101010;
         rom[429] = 24'b111111100111001001110100;
         rom[430] = 24'b111111011011010000011110;
         rom[431] = 24'b111111101110101010001101;
         rom[432] = 24'b111111110011011101101111;
         rom[433] = 24'b000000000011010001010110;
         rom[434] = 24'b111111111111010011111000;
         rom[435] = 24'b000000001101000101011111;
         rom[436] = 24'b000000001101110001001101;
         rom[437] = 24'b000000001100010111110010;
         rom[438] = 24'b000000011101010100011001;
         rom[439] = 24'b000000100110111000100010;
         rom[440] = 24'b000000100110110000001010;
         rom[441] = 24'b000000100010000110010001;
         rom[442] = 24'b000000100000000100001110;
         rom[443] = 24'b000000010010100100010000;
         rom[444] = 24'b000000100100101001110111;
         rom[445] = 24'b000000011001101010110110;
         rom[446] = 24'b000000001110000111000010;
         rom[447] = 24'b000000010011111111011001;
         rom[448] = 24'b000000001110011011010010;
         rom[449] = 24'b000000010100101000110101;
         rom[450] = 24'b111111110100011111111001;
         rom[451] = 24'b111111111101111110000011;
         rom[452] = 24'b111111110100010100010110;
         rom[453] = 24'b111111110000111100111101;
         rom[454] = 24'b111111101100101100000001;
         rom[455] = 24'b111111101101101000011100;
         rom[456] = 24'b111111010000011001010010;
         rom[457] = 24'b111111010010110101001010;
         rom[458] = 24'b111111010111010000001011;
         rom[459] = 24'b111111010000101001100110;
         rom[460] = 24'b111111001110101111110110;
         rom[461] = 24'b111111100010100110011010;
         rom[462] = 24'b111111101110011011011101;
         rom[463] = 24'b111111101011000100011000;
         rom[464] = 24'b111111011101111111010000;
         rom[465] = 24'b111111101101110011001001;
         rom[466] = 24'b111111111011001010101111;
         rom[467] = 24'b111111110110001100100111;
         rom[468] = 24'b000000010100010110111011;
         rom[469] = 24'b000000010010100110001000;
         rom[470] = 24'b000000010111001001010001;
         rom[471] = 24'b000000011000110100010000;
         rom[472] = 24'b000000100100110011110110;
         rom[473] = 24'b000000100100111100101101;
         rom[474] = 24'b000000011111010011111010;
         rom[475] = 24'b000000100010100100000111;
         rom[476] = 24'b000000110100001001010000;
         rom[477] = 24'b000000011010101011100111;
         rom[478] = 24'b000000100011111101101101;
         rom[479] = 24'b000000101000110110111001;
         rom[480] = 24'b000000010010011111100101;
         rom[481] = 24'b000000010101000111111001;
         rom[482] = 24'b000000011100011011010001;
         rom[483] = 24'b111111111001010101111100;
         rom[484] = 24'b111111110101110101001111;
         rom[485] = 24'b000000000000011111101010;
         rom[486] = 24'b111111111001010010100010;
         rom[487] = 24'b111111100110111100110110;
         rom[488] = 24'b111111100001101010000000;
         rom[489] = 24'b111111010011110100011000;
         rom[490] = 24'b111111100011011001000111;
         rom[491] = 24'b111111101000101101010100;
         rom[492] = 24'b111111011101011100000100;
         rom[493] = 24'b111111010110001110110111;
         rom[494] = 24'b111111011101101111000100;
         rom[495] = 24'b111111011100110000101101;
         rom[496] = 24'b111111100110110001101100;
         rom[497] = 24'b111111101100111000001000;
         rom[498] = 24'b111111110110111100000110;
         rom[499] = 24'b111111101100000001101110;
         rom[500] = 24'b000000001010000111000011;
         rom[501] = 24'b000000000101111001111000;
         rom[502] = 24'b000000001000011101101011;
         rom[503] = 24'b000000010101001111000000;
         rom[504] = 24'b000000010011001111100001;
         rom[505] = 24'b000000011001010010110000;
         rom[506] = 24'b000000011101101101111101;
         rom[507] = 24'b000000011000000100010100;
         rom[508] = 24'b000000100000111010001011;
         rom[509] = 24'b000000101011111001111110;
         rom[510] = 24'b000000101110110010000011;
         rom[511] = 24'b000000100000000101010100;
         rom[512] = 24'b000000100001001111100010;
         rom[513] = 24'b000000010111001001011001;
         rom[514] = 24'b000000000101010001110101;
         rom[515] = 24'b000000001010100100011000;
         rom[516] = 24'b000000001111001101101100;
         rom[517] = 24'b111111111111110110001110;
         rom[518] = 24'b111111111010010011101101;
         rom[519] = 24'b111111101001111111000101;
         rom[520] = 24'b111111011110011010111000;
         rom[521] = 24'b111111100101000110001100;
         rom[522] = 24'b111111011111010101100111;
         rom[523] = 24'b111111010010011100111000;
         rom[524] = 24'b111111001111100100110000;
         rom[525] = 24'b111111010110111000000011;
         rom[526] = 24'b111111011110110011101000;
         rom[527] = 24'b111111100000011000101110;
         rom[528] = 24'b111111101000111011000000;
         rom[529] = 24'b111111011101011110110100;
         rom[530] = 24'b111111101001011110110111;
         rom[531] = 24'b111111100101001110110000;
         rom[532] = 24'b111111110100110100101010;
         rom[533] = 24'b111111110000100111111010;
         rom[534] = 24'b000000001111011110111010;
         rom[535] = 24'b000000001000010001001100;
         rom[536] = 24'b000000001111011111010110;
         rom[537] = 24'b000000011101010100011101;
         rom[538] = 24'b000000010111010110101000;
         rom[539] = 24'b000000011110100101010101;
         rom[540] = 24'b000000100000101001010010;
         rom[541] = 24'b000000100101010010000111;
         rom[542] = 24'b000000100011001001010111;
         rom[543] = 24'b000000110011011000111000;
         rom[544] = 24'b000000011111101100110001;
         rom[545] = 24'b000000011111011001101000;
         rom[546] = 24'b000000011101110100010010;
         rom[547] = 24'b000000010001110110101010;
         rom[548] = 24'b000000011000000000100110;
         rom[549] = 24'b000000000010111010001001;
         rom[550] = 24'b111111101110110001011100;
         rom[551] = 24'b111111111010000001011101;
         rom[552] = 24'b111111101111110000010010;
         rom[553] = 24'b111111101011100111101110;
         rom[554] = 24'b111111110101001110100000;
         rom[555] = 24'b111111101000010110001000;
         rom[556] = 24'b111111011111011110111011;
         rom[557] = 24'b111111100111011111110010;
         rom[558] = 24'b111111011000011011011100;
         rom[559] = 24'b111111011101100011111100;
         rom[560] = 24'b111111011100011111011101;
         rom[561] = 24'b111111110001001000000100;
         rom[562] = 24'b111111101000010010011011;
         rom[563] = 24'b111111101001110110011000;
         rom[564] = 24'b111111100011110001110111;
         rom[565] = 24'b111111110010100011101001;
         rom[566] = 24'b111111110010010011011000;
         rom[567] = 24'b000000001001011100000101;
         rom[568] = 24'b000000000110001101101111;
         rom[569] = 24'b000000000010000110001111;
         rom[570] = 24'b000000001101110101110010;
         rom[571] = 24'b000000011110001010100010;
         rom[572] = 24'b000000011001111101111001;
         rom[573] = 24'b000000100100100010101010;
         rom[574] = 24'b000000110001111101111100;
         rom[575] = 24'b000000101011011011110101;
         rom[576] = 24'b000000110010001111101010;
         rom[577] = 24'b000000011101111000011000;
         rom[578] = 24'b000000100001110101011101;
         rom[579] = 24'b000000010011111010110010;
         rom[580] = 24'b000000010100011110010010;
         rom[581] = 24'b000000010000101100101011;
         rom[582] = 24'b000000000110110101110011;
         rom[583] = 24'b000000001011111001001000;
         rom[584] = 24'b000000000111001100001100;
         rom[585] = 24'b111111110111001010101000;
         rom[586] = 24'b111111101011011010101101;
         rom[587] = 24'b111111100111101001111100;
         rom[588] = 24'b111111011100110011010000;
         rom[589] = 24'b111111011101100101101000;
         rom[590] = 24'b111111011010100111110001;
         rom[591] = 24'b111111100101011001101001;
         rom[592] = 24'b111111010111111110101111;
         rom[593] = 24'b111111011010000010001110;
         rom[594] = 24'b111111101010010000100011;
         rom[595] = 24'b111111010111100110111001;
         rom[596] = 24'b111111100100010000111010;
         rom[597] = 24'b111111101110011011010111;
         rom[598] = 24'b111111101101111101101110;
         rom[599] = 24'b000000000010000000111000;
         rom[600] = 24'b111111111001110110110110;
         rom[601] = 24'b000000000100011100011010;
         rom[602] = 24'b111111111111100010101110;
         rom[603] = 24'b000000010010011000110100;
         rom[604] = 24'b000000100011100010010011;
         rom[605] = 24'b000000011011101001110001;
         rom[606] = 24'b000000101111000001000001;
         rom[607] = 24'b000000100010010100111101;
         rom[608] = 24'b000000010110101011010000;
         rom[609] = 24'b000000100101010111000001;
         rom[610] = 24'b000000100111111101010101;
         rom[611] = 24'b000000100000011001101101;
         rom[612] = 24'b000000011011111010011010;
         rom[613] = 24'b000000010110001101111100;
         rom[614] = 24'b000000011101011011110000;
         rom[615] = 24'b000000001100001000001010;
         rom[616] = 24'b000000000100001011111010;
         rom[617] = 24'b000000001011101001101011;
         rom[618] = 24'b111111101111100011111000;
         rom[619] = 24'b111111100100100000000100;
         rom[620] = 24'b111111110000010111001001;
         rom[621] = 24'b111111100101100101001100;
         rom[622] = 24'b111111100011011000110011;
         rom[623] = 24'b111111011111010000111100;
         rom[624] = 24'b111111011011010011001110;
         rom[625] = 24'b111111011010110010001110;
         rom[626] = 24'b111111001100000100010110;
         rom[627] = 24'b111111010010110010011010;
         rom[628] = 24'b111111100100110100001101;
         rom[629] = 24'b111111110000000000100111;
         rom[630] = 24'b111111100001010000100110;
         rom[631] = 24'b111111100101010010101001;
         rom[632] = 24'b111111111110110011101111;
         rom[633] = 24'b111111111101101100011010;
         rom[634] = 24'b000000000001110100001101;
         rom[635] = 24'b000000001011111011100000;
         rom[636] = 24'b000000011000100010010111;
         rom[637] = 24'b000000010101110101110100;
         rom[638] = 24'b000000010011111011100010;
         rom[639] = 24'b000000101100011001001011;
         rom[640] = 24'b000000011110011001001110;
         rom[641] = 24'b000000011010111111000011;
         rom[642] = 24'b000000100001100110011101;
         rom[643] = 24'b000000101000101101001101;
         rom[644] = 24'b000000011001110011010111;
         rom[645] = 24'b000000011101100110001100;
         rom[646] = 24'b000000011001011111000000;
         rom[647] = 24'b000000010110001101010010;
         rom[648] = 24'b000000000110111001011101;
         rom[649] = 24'b000000000011010101110111;
         rom[650] = 24'b111111111001110110100000;
         rom[651] = 24'b111111111001101000101001;
         rom[652] = 24'b111111111111010100000111;
         rom[653] = 24'b111111110100000001101001;
         rom[654] = 24'b111111111000101000110100;
         rom[655] = 24'b111111100010110101000001;
         rom[656] = 24'b111111011111101111010101;
         rom[657] = 24'b111111011001100010010100;
         rom[658] = 24'b111111011000101110111111;
         rom[659] = 24'b111111011100000001011100;
         rom[660] = 24'b111111011110000011000101;
         rom[661] = 24'b111111011011000111100001;
         rom[662] = 24'b111111100101101111000111;
         rom[663] = 24'b111111101011101010110100;
         rom[664] = 24'b111111110000111101001110;
         rom[665] = 24'b111111110100000111010000;
         rom[666] = 24'b000000000011001101000000;
         rom[667] = 24'b000000000010000011011001;
         rom[668] = 24'b000000001000011011000100;
         rom[669] = 24'b000000000011101011000011;
         rom[670] = 24'b000000010011001011111011;
         rom[671] = 24'b000000101010000111110100;
         rom[672] = 24'b000000100111000011100010;
         rom[673] = 24'b000000010001101001100001;
         rom[674] = 24'b000000101101010001101011;
         rom[675] = 24'b000000101001101000100010;
         rom[676] = 24'b000000011011111101111110;
         rom[677] = 24'b000000100011011101011011;
         rom[678] = 24'b000000100000111101001010;
         rom[679] = 24'b000000100110110101101111;
         rom[680] = 24'b000000010001000111010101;
         rom[681] = 24'b000000000111100111010111;
         rom[682] = 24'b000000001101100110110111;
         rom[683] = 24'b000000001000101100111101;
         rom[684] = 24'b111111110111110000111111;
         rom[685] = 24'b111111111110010010101101;
         rom[686] = 24'b111111101011110000101010;
         rom[687] = 24'b111111100111001100010011;
         rom[688] = 24'b111111011010000100100001;
         rom[689] = 24'b111111100111100010100111;
         rom[690] = 24'b111111100100000001011101;
         rom[691] = 24'b111111011100111001110111;
         rom[692] = 24'b111111001101010011100011;
         rom[693] = 24'b111111100100111000010111;
         rom[694] = 24'b111111100100010111110000;
         rom[695] = 24'b111111100000101001010111;
         rom[696] = 24'b111111100001111100001100;
         rom[697] = 24'b111111100110010010011100;
         rom[698] = 24'b111111100111010011110100;
         rom[699] = 24'b111111101011100101110011;
         rom[700] = 24'b111111111111100110101011;
         rom[701] = 24'b000000000000101011010110;
         rom[702] = 24'b000000010000010011111001;
         rom[703] = 24'b000000010110111110100001;
         rom[704] = 24'b000000010110011001010100;
         rom[705] = 24'b000000011110111100100001;
         rom[706] = 24'b000000100110111101111101;
         rom[707] = 24'b000000100100101100111000;
         rom[708] = 24'b000000101101100000000001;
         rom[709] = 24'b000000100100100101110100;
         rom[710] = 24'b000000011110100100100111;
         rom[711] = 24'b000000010111111011000000;
         rom[712] = 24'b000000010001000110101011;
         rom[713] = 24'b000000011100011101100100;
         rom[714] = 24'b000000011010111110111001;
         rom[715] = 24'b000000010110110110000111;
         rom[716] = 24'b111111111111100100110110;
         rom[717] = 24'b000000000010111011100001;
         rom[718] = 24'b111111101111101111101011;
         rom[719] = 24'b111111110110111111100011;
         rom[720] = 24'b111111100111110100101011;
         rom[721] = 24'b111111110100100110000110;
         rom[722] = 24'b111111100110011011101111;
         rom[723] = 24'b111111011001100110110011;
         rom[724] = 24'b111111101000100101100101;
         rom[725] = 24'b111111100000001010111010;
         rom[726] = 24'b111111100110000010011111;
         rom[727] = 24'b111111011010010011110001;
         rom[728] = 24'b111111101001101101100011;
         rom[729] = 24'b111111110001111111010001;
         rom[730] = 24'b111111100110100010000110;
         rom[731] = 24'b111111101010101000011011;
         rom[732] = 24'b111111111111101100010111;
         rom[733] = 24'b111111111001010011001011;
         rom[734] = 24'b000000000111010000000101;
         rom[735] = 24'b000000000111000000000000;
         rom[736] = 24'b000000010011010110010100;
         rom[737] = 24'b000000011011010101100111;
         rom[738] = 24'b000000100000111001110100;
         rom[739] = 24'b000000010010000000100001;
         rom[740] = 24'b000000011000100010101100;
         rom[741] = 24'b000000011010100111110000;
         rom[742] = 24'b000000101001101010011110;
         rom[743] = 24'b000000101001000111100011;
         rom[744] = 24'b000000011101011110011101;
         rom[745] = 24'b000000100010000111001100;
         rom[746] = 24'b000000100011010010100100;
         rom[747] = 24'b000000010010000111100010;
         rom[748] = 24'b000000001101000011010101;
         rom[749] = 24'b000000000101110010001011;
         rom[750] = 24'b111111110110010010111111;
         rom[751] = 24'b111111111100101101000000;
         rom[752] = 24'b111111100010011100101011;
         rom[753] = 24'b111111110111010101110000;
         rom[754] = 24'b111111110010101111011010;
         rom[755] = 24'b111111100111110101110111;
         rom[756] = 24'b111111100100100011111011;
         rom[757] = 24'b111111011110110011111111;
         rom[758] = 24'b111111101101011111011000;
         rom[759] = 24'b111111011001101110100001;
         rom[760] = 24'b111111010100010000100010;
         rom[761] = 24'b111111101011111001111110;
         rom[762] = 24'b111111011110110000001100;
         rom[763] = 24'b111111101111010110000011;
         rom[764] = 24'b111111100011101011001000;
         rom[765] = 24'b111111101011111100100000;
         rom[766] = 24'b000000000010110010010011;
         rom[767] = 24'b000000000001001011101010;
         rom[768] = 24'b000000001111101001110111;
         rom[769] = 24'b000000010000011010011000;
         rom[770] = 24'b000000011110001010100110;
         rom[771] = 24'b000000101001010111010111;
         rom[772] = 24'b000000010110111011010101;
         rom[773] = 24'b000000101000000100110100;
         rom[774] = 24'b000000011111111011100000;
         rom[775] = 24'b000000100111011100110111;
         rom[776] = 24'b000000100001101110001101;
         rom[777] = 24'b000000100101100000000101;
         rom[778] = 24'b000000100001110001000001;
         rom[779] = 24'b000000011101010000011010;
         rom[780] = 24'b000000001011101010110100;
         rom[781] = 24'b000000000100010100100000;
         rom[782] = 24'b000000010001011010101010;
         rom[783] = 24'b000000000100100000001000;
         rom[784] = 24'b111111111000010101111001;
         rom[785] = 24'b000000000011101100101011;
         rom[786] = 24'b111111110011001100010101;
         rom[787] = 24'b111111110101010011000100;
         rom[788] = 24'b111111100101101011000101;
         rom[789] = 24'b111111011111100000110001;
         rom[790] = 24'b111111011101011111110010;
         rom[791] = 24'b111111010010111110001100;
         rom[792] = 24'b111111100000111010111101;
         rom[793] = 24'b111111011100110111101000;
         rom[794] = 24'b111111011111100010001000;
         rom[795] = 24'b111111110001011000011011;
         rom[796] = 24'b111111110010010000001000;
         rom[797] = 24'b111111110000011101110011;
         rom[798] = 24'b111111110100000000101101;
         rom[799] = 24'b000000000110000110100011;
         rom[800] = 24'b111111111011011000101001;
         rom[801] = 24'b000000001001010011011110;
         rom[802] = 24'b000000000100111101100001;
         rom[803] = 24'b000000011110001100101110;
         rom[804] = 24'b000000100010111100100110;
         rom[805] = 24'b000000011001101100000010;
         rom[806] = 24'b000000011010110000010101;
         rom[807] = 24'b000000100111111100001110;
         rom[808] = 24'b000000101100000010010101;
         rom[809] = 24'b000000100000101001101101;
         rom[810] = 24'b000000010110001001110101;
         rom[811] = 24'b000000100001010110100101;
         rom[812] = 24'b000000011000101101010000;
         rom[813] = 24'b000000010010000110010000;
         rom[814] = 24'b000000001011110000100011;
         rom[815] = 24'b000000001111010100001100;
         rom[816] = 24'b000000001010000101000001;
         rom[817] = 24'b111111111001010001100100;
         rom[818] = 24'b111111101100110000010111;
         rom[819] = 24'b111111101010110011010101;
         rom[820] = 24'b111111101110001100011011;
         rom[821] = 24'b111111100000011111000110;
         rom[822] = 24'b111111101010001001011011;
         rom[823] = 24'b111111011101100101101111;
         rom[824] = 24'b111111100001000101110111;
         rom[825] = 24'b111111011011010000100000;
         rom[826] = 24'b111111011111110001001000;
         rom[827] = 24'b111111010001101001001110;
         rom[828] = 24'b111111101001001011011111;
         rom[829] = 24'b111111100101111100000000;
         rom[830] = 24'b111111101111101100100010;
         rom[831] = 24'b111111101000001111000010;
         rom[832] = 24'b111111111100101101111010;
         rom[833] = 24'b000000000100001011101000;
         rom[834] = 24'b111111111101100000111100;
         rom[835] = 24'b000000001001110000010010;
         rom[836] = 24'b000000010001011010000110;
         rom[837] = 24'b000000010100100101000101;
         rom[838] = 24'b000000100111000110100110;
         rom[839] = 24'b000000100001011011010011;
         rom[840] = 24'b000000101000011001100110;
         rom[841] = 24'b000000100001001110101111;
         rom[842] = 24'b000000110001000111010010;
         rom[843] = 24'b000000100110010000001010;
         rom[844] = 24'b000000100001100101000101;
         rom[845] = 24'b000000011110001101000000;
         rom[846] = 24'b000000011011000111001101;
         rom[847] = 24'b000000001001100000100111;
         rom[848] = 24'b000000010010101100111011;
         rom[849] = 24'b111111111111010010001110;
         rom[850] = 24'b000000000000100001001000;
         rom[851] = 24'b111111111110011011011110;
         rom[852] = 24'b111111101110000000110010;
         rom[853] = 24'b111111101010111101011010;
         rom[854] = 24'b111111011111000000011001;
         rom[855] = 24'b111111100011110011111010;
         rom[856] = 24'b111111100111000000010101;
         rom[857] = 24'b111111100001111101110111;
         rom[858] = 24'b111111010111010000000010;
         rom[859] = 24'b111111011011101001100010;
         rom[860] = 24'b111111011010101111000000;
         rom[861] = 24'b111111011010000101111110;
         rom[862] = 24'b111111100110011101110000;
         rom[863] = 24'b111111110001111101000010;
         rom[864] = 24'b111111101101100101110101;
         rom[865] = 24'b111111101101111000110001;
         rom[866] = 24'b111111111110010111111010;
         rom[867] = 24'b000000000101011110001111;
         rom[868] = 24'b000000001110010100001110;
         rom[869] = 24'b000000001001100010000110;
         rom[870] = 24'b000000010110001000000011;
         rom[871] = 24'b000000010010110001110011;
         rom[872] = 24'b000000100111000101110101;
         rom[873] = 24'b000000011001011011001000;
         rom[874] = 24'b000000011111010110101100;
         rom[875] = 24'b000000011111101111101001;
         rom[876] = 24'b000000100100100010011111;
         rom[877] = 24'b000000101000000111110100;
         rom[878] = 24'b000000010111111100100110;
         rom[879] = 24'b000000100100111110011001;
         rom[880] = 24'b000000001010101111101111;
         rom[881] = 24'b000000010001001010000010;
         rom[882] = 24'b000000001011111111101101;
         rom[883] = 24'b000000000100011010001111;
         rom[884] = 24'b111111111100100001111000;
         rom[885] = 24'b111111110101100110101111;
         rom[886] = 24'b111111110000010110010001;
         rom[887] = 24'b111111101000101000011011;
         rom[888] = 24'b111111011110100101110101;
         rom[889] = 24'b111111100110110011000101;
         rom[890] = 24'b111111010111101100000101;
         rom[891] = 24'b111111100001111101111010;
         rom[892] = 24'b111111011101110101101011;
         rom[893] = 24'b111111100011111001001010;
         rom[894] = 24'b111111011000011101001100;
         rom[895] = 24'b111111100111110111101000;
         rom[896] = 24'b111111011010100000111110;
         rom[897] = 24'b111111101001100001000110;
         rom[898] = 24'b111111111011000110000010;
         rom[899] = 24'b000000000111000011000000;
         rom[900] = 24'b111111111110010101001001;
         rom[901] = 24'b000000000101000100000010;
         rom[902] = 24'b000000010000101101011110;
         rom[903] = 24'b000000001011111010100100;
         rom[904] = 24'b000000001011001001010001;
         rom[905] = 24'b000000100010111001010010;
         rom[906] = 24'b000000011100111010000110;
         rom[907] = 24'b000000011001010001101110;
         rom[908] = 24'b000000100100010000010110;
         rom[909] = 24'b000000100110011000111100;
         rom[910] = 24'b000000011011001010011100;
         rom[911] = 24'b000000010110110110110001;
         rom[912] = 24'b000000100010010001011000;
         rom[913] = 24'b000000011110101001110101;
         rom[914] = 24'b000000001010001010001000;
         rom[915] = 24'b000000010011110110001011;
         rom[916] = 24'b000000000011011001111001;
         rom[917] = 24'b000000000111101001000000;
         rom[918] = 24'b111111111100101101101001;
         rom[919] = 24'b111111110110111011011110;
         rom[920] = 24'b111111101100100111100101;
         rom[921] = 24'b111111011010100100110111;
         rom[922] = 24'b111111100101000011001110;
         rom[923] = 24'b111111100110111101101000;
         rom[924] = 24'b111111011101011001100110;
         rom[925] = 24'b111111011001010101110100;
         rom[926] = 24'b111111101101101000111011;
         rom[927] = 24'b111111011110001100111000;
         rom[928] = 24'b111111011110010010011111;
         rom[929] = 24'b111111101000011100110001;
         rom[930] = 24'b111111100101000000001100;
         rom[931] = 24'b111111110011011001111000;
         rom[932] = 24'b111111101111010101000000;
         rom[933] = 24'b111111111110010110011000;
         rom[934] = 24'b000000001110011110111010;
         rom[935] = 24'b000000010011010010001001;
         rom[936] = 24'b000000001101000010110111;
         rom[937] = 24'b000000010100100111111111;
         rom[938] = 24'b000000011110100011111001;
         rom[939] = 24'b000000100001110100010110;
         rom[940] = 24'b000000011100011111000101;
         rom[941] = 24'b000000100010001001110010;
         rom[942] = 24'b000000100010000100110111;
         rom[943] = 24'b000000100000001000010110;
         rom[944] = 24'b000000011111110110100011;
         rom[945] = 24'b000000011101011010100010;
         rom[946] = 24'b000000010011101111101011;
         rom[947] = 24'b000000001011101010110101;
         rom[948] = 24'b000000001100100010110101;
         rom[949] = 24'b000000010000111100111001;
         rom[950] = 24'b111111111011110000110100;
         rom[951] = 24'b111111110101110011001001;
         rom[952] = 24'b111111101011101000011001;
         rom[953] = 24'b111111101001111010010011;
         rom[954] = 24'b111111101010011111100011;
         rom[955] = 24'b111111100001000010111110;
         rom[956] = 24'b111111100010110101101001;
         rom[957] = 24'b111111100111011100101001;
         rom[958] = 24'b111111011110011101110000;
         rom[959] = 24'b111111100011010010010010;
         rom[960] = 24'b111111101000101011100110;
         rom[961] = 24'b111111011110000101001011;
         rom[962] = 24'b111111011100001000010110;
         rom[963] = 24'b111111110011101101101110;
         rom[964] = 24'b111111110110101001011011;
         rom[965] = 24'b111111111011100010010100;
         rom[966] = 24'b000000000101111011010110;
         rom[967] = 24'b111111110111011111111110;
         rom[968] = 24'b111111111111010111111011;
         rom[969] = 24'b000000010100000001110010;
         rom[970] = 24'b000000001011111100011011;
         rom[971] = 24'b000000100111000010110000;
         rom[972] = 24'b000000100110001101010010;
         rom[973] = 24'b000000101100011100100000;
         rom[974] = 24'b000000011000110111001001;
         rom[975] = 24'b000000100010010011101110;
         rom[976] = 24'b000000101100010010111001;
         rom[977] = 24'b000000100000100000010001;
         rom[978] = 24'b000000011110001100011011;
         rom[979] = 24'b000000010001010000011101;
         rom[980] = 24'b000000001111100100001011;
         rom[981] = 24'b000000010101001011101101;
         rom[982] = 24'b000000001100110011110101;
         rom[983] = 24'b111111111111101110010100;
         rom[984] = 24'b111111111101111110101000;
         rom[985] = 24'b111111110111110100101011;
         rom[986] = 24'b111111101101101011101111;
         rom[987] = 24'b111111100111000010010011;
         rom[988] = 24'b111111011000110101010001;
         rom[989] = 24'b111111010000111010011010;
         rom[990] = 24'b111111011100100010101000;
         rom[991] = 24'b111111100001001011000001;
         rom[992] = 24'b111111010000000010000000;
         rom[993] = 24'b111111001111110000001001;
         rom[994] = 24'b111111011001110110100011;
         rom[995] = 24'b111111011011100101101010;
         rom[996] = 24'b111111110001011110110111;
         rom[997] = 24'b111111100101011110100001;
         rom[998] = 24'b111111111110010011110101;
         rom[999] = 24'b000000000111111010101000;
         rom[1000] = 24'b000000001011110100011110;
         rom[1001] = 24'b000000010011101011000000;
         rom[1002] = 24'b000000000001111101000110;
         rom[1003] = 24'b000000000111100001001010;
         rom[1004] = 24'b000000010010010100111111;
         rom[1005] = 24'b000000010101001001001010;
         rom[1006] = 24'b000000100001100000111001;
         rom[1007] = 24'b000000100010011101000011;
         rom[1008] = 24'b000000100100011100010011;
         rom[1009] = 24'b000000100111101010111100;
         rom[1010] = 24'b000000010111000100000000;
         rom[1011] = 24'b000000011011001010111001;
         rom[1012] = 24'b000000100000110000110010;
         rom[1013] = 24'b000000011110111100010010;
         rom[1014] = 24'b000000011001000001000110;
         rom[1015] = 24'b000000010000110011001101;
         rom[1016] = 24'b000000010001000010100111;
         rom[1017] = 24'b000000001001010011000100;
         rom[1018] = 24'b111111101111100110101011;
         rom[1019] = 24'b111111101111011011110111;
         rom[1020] = 24'b111111100101101001100001;
         rom[1021] = 24'b111111011000001110100000;
         rom[1022] = 24'b111111011010000010001011;
         rom[1023] = 24'b111111011000000010101111;
         rom[1024] = 24'b111111010101110111000110;
         rom[1025] = 24'b111111100000000100000001;
         rom[1026] = 24'b111111100011101111100011;
         rom[1027] = 24'b111111101100011100001100;
         rom[1028] = 24'b111111101011100110001010;
         rom[1029] = 24'b111111101011010011111010;
         rom[1030] = 24'b111111110100100111011011;
         rom[1031] = 24'b111111100111101111110011;
         rom[1032] = 24'b111111110010101000001001;
         rom[1033] = 24'b111111111111011000001001;
         rom[1034] = 24'b111111111100001000111010;
         rom[1035] = 24'b000000010010010010001011;
         rom[1036] = 24'b000000001100110111100100;
         rom[1037] = 24'b000000011110001100011100;
         rom[1038] = 24'b000000011001111011001000;
         rom[1039] = 24'b000000100111011110100110;
         rom[1040] = 24'b000000100000010001010111;
         rom[1041] = 24'b000000100101111001111111;
         rom[1042] = 24'b000000100110111000011001;
         rom[1043] = 24'b000000101010001000011010;
         rom[1044] = 24'b000000101001001001100001;
         rom[1045] = 24'b000000011011101011101000;
         rom[1046] = 24'b000000011010111001000111;
         rom[1047] = 24'b000000010110101110011000;
         rom[1048] = 24'b000000001111011100110101;
         rom[1049] = 24'b000000001000100001110010;
         rom[1050] = 24'b111111111110111010000101;
         rom[1051] = 24'b111111110100010100011000;
         rom[1052] = 24'b111111110100011101001011;
         rom[1053] = 24'b111111101001010011010100;
         rom[1054] = 24'b111111101001100110100101;
         rom[1055] = 24'b111111110001010101111001;
         rom[1056] = 24'b111111100011100101000001;
         rom[1057] = 24'b111111100110100001001110;
         rom[1058] = 24'b111111101000010001010111;
         rom[1059] = 24'b111111010111101100111001;
         rom[1060] = 24'b111111100001011110001111;
         rom[1061] = 24'b111111100000100101101000;
         rom[1062] = 24'b111111101110001111000001;
         rom[1063] = 24'b111111110011001101111100;
         rom[1064] = 24'b111111101101111110010011;
         rom[1065] = 24'b111111110100101111011000;
         rom[1066] = 24'b111111110010000000001000;
         rom[1067] = 24'b111111111010101001000001;
         rom[1068] = 24'b000000000100011010001110;
         rom[1069] = 24'b000000001011001010100010;
         rom[1070] = 24'b000000011001000100101000;
         rom[1071] = 24'b000000011000010010000010;
         rom[1072] = 24'b000000011001011011000011;
         rom[1073] = 24'b000000100000000001011000;
         rom[1074] = 24'b000000100101100001000011;
         rom[1075] = 24'b000000100100110000000010;
         rom[1076] = 24'b000000101000010110111110;
         rom[1077] = 24'b000000100001111001011101;
         rom[1078] = 24'b000000011111011010010010;
         rom[1079] = 24'b000000100100101000001011;
         rom[1080] = 24'b000000001110001110101101;
         rom[1081] = 24'b000000010111010111010101;
         rom[1082] = 24'b000000011101000001001010;
         rom[1083] = 24'b111111111101011111100100;
         rom[1084] = 24'b000000010000010011001111;
         rom[1085] = 24'b111111111011110110001111;
         rom[1086] = 24'b111111100010110001101100;
         rom[1087] = 24'b111111010100101011100010;
         rom[1088] = 24'b111111100000100001111011;
         rom[1089] = 24'b111111010011001101011110;
         rom[1090] = 24'b111111100100111011110011;
         rom[1091] = 24'b111111010100100110001110;
         rom[1092] = 24'b111111100110100110010110;
         rom[1093] = 24'b111111101000001010001110;
         rom[1094] = 24'b111111011001000100010100;
         rom[1095] = 24'b111111100000110000000010;
         rom[1096] = 24'b111111010101000110000010;
         rom[1097] = 24'b111111110000111111111101;
         rom[1098] = 24'b111111110100110110010010;
         rom[1099] = 24'b111111110101101000011001;
         rom[1100] = 24'b111111111000011010100110;
         rom[1101] = 24'b000000001101100110010001;
         rom[1102] = 24'b000000010000101110011001;
         rom[1103] = 24'b000000011100100110011110;
         rom[1104] = 24'b000000010101110101011001;
         rom[1105] = 24'b000000100000100110100100;
         rom[1106] = 24'b000000101001101101011101;
         rom[1107] = 24'b000000011101100110101101;
         rom[1108] = 24'b000000100010111011011111;
         rom[1109] = 24'b000000100010101100101011;
         rom[1110] = 24'b000000101010010001110010;
         rom[1111] = 24'b000000011111001111001000;
         rom[1112] = 24'b000000010001111110111101;
         rom[1113] = 24'b000000010001010010000100;
         rom[1114] = 24'b000000010110111110010001;
         rom[1115] = 24'b000000010011101111101000;
         rom[1116] = 24'b111111111111011001100111;
         rom[1117] = 24'b111111111101100001101010;
         rom[1118] = 24'b111111110010010110101100;
         rom[1119] = 24'b111111110011101011010111;
         rom[1120] = 24'b111111110111010010000011;
         rom[1121] = 24'b111111101111010011000001;
         rom[1122] = 24'b111111100100011001011101;
         rom[1123] = 24'b111111010110111101100100;
         rom[1124] = 24'b111111010101110010001010;
         rom[1125] = 24'b111111010111000010011011;
         rom[1126] = 24'b111111010001111110001000;
         rom[1127] = 24'b111111011010110001001110;
         rom[1128] = 24'b111111101000000101101111;
         rom[1129] = 24'b111111011010111011011011;
         rom[1130] = 24'b111111101111011001000010;
         rom[1131] = 24'b111111101010010011101010;
         rom[1132] = 24'b111111110100010111000100;
         rom[1133] = 24'b111111111001011000010111;
         rom[1134] = 24'b111111111000000000100001;
         rom[1135] = 24'b000000001110011000000111;
         rom[1136] = 24'b000000001110100011001000;
         rom[1137] = 24'b000000001001011001011110;
         rom[1138] = 24'b000000011111000110111110;
         rom[1139] = 24'b000000100101111000110000;
         rom[1140] = 24'b000000110011011000001000;
         rom[1141] = 24'b000000011111001111010001;
         rom[1142] = 24'b000000100000110100101011;
         rom[1143] = 24'b000000100101000000000100;
         rom[1144] = 24'b000000011110010101000011;
         rom[1145] = 24'b000000011111000000010011;
         rom[1146] = 24'b000000011011101110010011;
         rom[1147] = 24'b000000010100111101011111;
         rom[1148] = 24'b000000011110111001100110;
         rom[1149] = 24'b111111111110011010001101;
         rom[1150] = 24'b111111111111011001001011;
         rom[1151] = 24'b111111111010011010100011;
         rom[1152] = 24'b111111101100011101000101;
         rom[1153] = 24'b111111111101001111101110;
         rom[1154] = 24'b111111100100111101001000;
         rom[1155] = 24'b111111011100111010110011;
         rom[1156] = 24'b111111010010001110101010;
         rom[1157] = 24'b111111100000000111110101;
         rom[1158] = 24'b111111011101011001011110;
         rom[1159] = 24'b111111011000001111101010;
         rom[1160] = 24'b111111100100011101011100;
         rom[1161] = 24'b111111101000101110110010;
         rom[1162] = 24'b111111100111110110111100;
         rom[1163] = 24'b111111100010101001011000;
         rom[1164] = 24'b111111101010111011111100;
         rom[1165] = 24'b111111110001111100111111;
         rom[1166] = 24'b000000000101110100110010;
         rom[1167] = 24'b000000001100100010101010;
         rom[1168] = 24'b000000010010101011101010;
         rom[1169] = 24'b000000011011101011101110;
         rom[1170] = 24'b000000001101110010101010;
         rom[1171] = 24'b000000011010100101011000;
         rom[1172] = 24'b000000010010111110001101;
         rom[1173] = 24'b000000101101010000111011;
         rom[1174] = 24'b000000100010100000000000;
         rom[1175] = 24'b000000100101011000101011;
         rom[1176] = 24'b000000101010000101000110;
         rom[1177] = 24'b000000011101000001001111;
         rom[1178] = 24'b000000011101111101001101;
         rom[1179] = 24'b000000011010111100010110;
         rom[1180] = 24'b000000010111000000011100;
         rom[1181] = 24'b000000001110111000100001;
         rom[1182] = 24'b000000001011000101110101;
         rom[1183] = 24'b000000000001110111000011;
         rom[1184] = 24'b111111111100010011011100;
         rom[1185] = 24'b111111111001100110000100;
         rom[1186] = 24'b111111101101011010110000;
         rom[1187] = 24'b111111100000000111010101;
         rom[1188] = 24'b111111100101001011001101;
         rom[1189] = 24'b111111100000110000110010;
         rom[1190] = 24'b111111010100110010010001;
         rom[1191] = 24'b111111011000110000101010;
         rom[1192] = 24'b111111100010100000101100;
         rom[1193] = 24'b111111010110010110001000;
         rom[1194] = 24'b111111011101010101110101;
         rom[1195] = 24'b111111011110011110011011;
         rom[1196] = 24'b111111011101011010000011;
         rom[1197] = 24'b111111100010011001011000;
         rom[1198] = 24'b111111110010001110110000;
         rom[1199] = 24'b111111110111101100100001;
         rom[1200] = 24'b111111111101101010010011;
         rom[1201] = 24'b000000001111011111111111;
         rom[1202] = 24'b000000010011001000000101;
         rom[1203] = 24'b000000011101101101001001;
         rom[1204] = 24'b000000100001000110110101;
         rom[1205] = 24'b000000100101000011000010;
         rom[1206] = 24'b000000011101111111110001;
         rom[1207] = 24'b000000100001111101110001;
         rom[1208] = 24'b000000011010110000100110;
         rom[1209] = 24'b000000100101011101011001;
         rom[1210] = 24'b000000011101000010001100;
         rom[1211] = 24'b000000100010010011110011;
         rom[1212] = 24'b000000011101000110110010;
         rom[1213] = 24'b000000100111010001001011;
         rom[1214] = 24'b000000011001010101001110;
         rom[1215] = 24'b000000001001000110011110;
         rom[1216] = 24'b111111111011011011001101;
         rom[1217] = 24'b111111110000101101000011;
         rom[1218] = 24'b111111111001000110011100;
         rom[1219] = 24'b111111111000101110001100;
         rom[1220] = 24'b111111101010011000010111;
         rom[1221] = 24'b111111011110000100000010;
         rom[1222] = 24'b111111010100011100011101;
         rom[1223] = 24'b111111010110000010000000;
         rom[1224] = 24'b111111011110000100001000;
         rom[1225] = 24'b111111011010000001000001;
         rom[1226] = 24'b111111011010001000000011;
         rom[1227] = 24'b111111101101001000000000;
         rom[1228] = 24'b111111100111111110110100;
         rom[1229] = 24'b111111101011100111101000;
         rom[1230] = 24'b111111100110001001011011;
         rom[1231] = 24'b111111111100110000110011;
         rom[1232] = 24'b000000000100101101000101;
         rom[1233] = 24'b111111111110110100101101;
         rom[1234] = 24'b000000000111110000010011;
         rom[1235] = 24'b000000000110001011111110;
         rom[1236] = 24'b000000010001001000011010;
         rom[1237] = 24'b000000011101011000000111;
         rom[1238] = 24'b000000011100001110000000;
         rom[1239] = 24'b000000100000111001100011;
         rom[1240] = 24'b000000101110011101001111;
         rom[1241] = 24'b000000011110111100000100;
         rom[1242] = 24'b000000011111001101000111;
         rom[1243] = 24'b000000101111010111110111;
         rom[1244] = 24'b000000100001010111100010;
         rom[1245] = 24'b000000011011011001110000;
         rom[1246] = 24'b000000010010011100110011;
         rom[1247] = 24'b000000011100000110110010;
         rom[1248] = 24'b000000010000000111111110;
         rom[1249] = 24'b000000000111011000000111;
         rom[1250] = 24'b111111111100101000011011;
         rom[1251] = 24'b111111110011011000001101;
         rom[1252] = 24'b111111101101100001101110;
         rom[1253] = 24'b111111101110011111111110;
         rom[1254] = 24'b111111101010011111001110;
         rom[1255] = 24'b111111011011101010110110;
         rom[1256] = 24'b111111011111011010101001;
         rom[1257] = 24'b111111010000110110011110;
         rom[1258] = 24'b111111010111000111000100;
         rom[1259] = 24'b111111011000001011100011;
         rom[1260] = 24'b111111010100001110111000;
         rom[1261] = 24'b111111100001001110000000;
         rom[1262] = 24'b111111011110010001101101;
         rom[1263] = 24'b111111100011110100111110;
         rom[1264] = 24'b111111101010110011010100;
         rom[1265] = 24'b111111110011110111000111;
         rom[1266] = 24'b111111110111011111000001;
         rom[1267] = 24'b000000000011110111111001;
         rom[1268] = 24'b111111111111111000001101;
         rom[1269] = 24'b000000011110011111111101;
         rom[1270] = 24'b000000011010101111010011;
         rom[1271] = 24'b000000001110001010010000;
         rom[1272] = 24'b000000011100110101001101;
         rom[1273] = 24'b000000100000001110100011;
         rom[1274] = 24'b000000101101100001101011;
         rom[1275] = 24'b000000100101111101001000;
         rom[1276] = 24'b000000101001000101000011;
         rom[1277] = 24'b000000011100110000011001;
         rom[1278] = 24'b000000011111110101011110;
         rom[1279] = 24'b000000011010000101000001;
         rom[1280] = 24'b000000010100111001011100;
         rom[1281] = 24'b000000010100110010100100;
         rom[1282] = 24'b111111111111100101110111;
         rom[1283] = 24'b000000000010000001111111;
         rom[1284] = 24'b000000001110000100110110;
         rom[1285] = 24'b111111110010011100101100;
         rom[1286] = 24'b111111111000101101011010;
         rom[1287] = 24'b111111101001001001000110;
         rom[1288] = 24'b111111011010110101100101;
         rom[1289] = 24'b111111011100011000001000;
         rom[1290] = 24'b111111011110100001100111;
         rom[1291] = 24'b111111010110010110001010;
         rom[1292] = 24'b111111011101100101101110;
         rom[1293] = 24'b111111100101011010111000;
         rom[1294] = 24'b111111100100111000100100;
         rom[1295] = 24'b111111011001010010010001;
         rom[1296] = 24'b111111101011001011000011;
         rom[1297] = 24'b111111111000011111011010;
         rom[1298] = 24'b111111110111110001000011;
         rom[1299] = 24'b111111111011111111000011;
         rom[1300] = 24'b111111110011111010001111;
         rom[1301] = 24'b000000000111111101111000;
         rom[1302] = 24'b000000100001001001010000;
         rom[1303] = 24'b000000101101001011110011;
         rom[1304] = 24'b000000110100101101111010;
         rom[1305] = 24'b000001000011101111111011;
         rom[1306] = 24'b000001000111110000100100;
         rom[1307] = 24'b000001011001000010010011;
         rom[1308] = 24'b000001010100010101101100;
         rom[1309] = 24'b000001101001101100010011;
         rom[1310] = 24'b000001101111000110100111;
         rom[1311] = 24'b000001101101110100111010;
         rom[1312] = 24'b000001111011010001010111;
         rom[1313] = 24'b000001101110100110001111;
         rom[1314] = 24'b000001111010010100011110;
         rom[1315] = 24'b000001111011111001010111;
         rom[1316] = 24'b000001111110001010101110;
         rom[1317] = 24'b000010000100001001000000;
         rom[1318] = 24'b000001111111000101010101;
         rom[1319] = 24'b000010000000010101001100;
         rom[1320] = 24'b000001111110101010010101;
         rom[1321] = 24'b000001110111000000001011;
         rom[1322] = 24'b000010000010010111011000;
         rom[1323] = 24'b000010000001001100011101;
         rom[1324] = 24'b000010001011010110011010;
         rom[1325] = 24'b000010010110111010000010;
         rom[1326] = 24'b000010010011111101010010;
         rom[1327] = 24'b000010100001000101110101;
         rom[1328] = 24'b000010100011100010110011;
         rom[1329] = 24'b000011000010010000101110;
         rom[1330] = 24'b000011001101001100100101;
         rom[1331] = 24'b000011010010100110001001;
         rom[1332] = 24'b000011011100000110010010;
         rom[1333] = 24'b000011101001100001001010;
         rom[1334] = 24'b000011111101010101010111;
         rom[1335] = 24'b000100001000010110110101;
         rom[1336] = 24'b000100000111100010100011;
         rom[1337] = 24'b000100101110000101110101;
         rom[1338] = 24'b000100110000011110110011;
         rom[1339] = 24'b000100110110011001101001;
         rom[1340] = 24'b000101001100110111111010;
         rom[1341] = 24'b000101001110101101101001;
         rom[1342] = 24'b000101001100101100000100;
         rom[1343] = 24'b000101011001110100110111;
         rom[1344] = 24'b000101100011011001000000;
         rom[1345] = 24'b000101100000010100111101;
         rom[1346] = 24'b000101110001100111001001;
         rom[1347] = 24'b000101101011011111001110;
         rom[1348] = 24'b000101101001011110101010;
         rom[1349] = 24'b000101101010100001110100;
         rom[1350] = 24'b000101111001011111110110;
         rom[1351] = 24'b000101100001100101010000;
         rom[1352] = 24'b000101110000011111010010;
         rom[1353] = 24'b000101111111111001111001;
         rom[1354] = 24'b000101101000100110000010;
         rom[1355] = 24'b000101110111000110011001;
         rom[1356] = 24'b000101110001101111001111;
         rom[1357] = 24'b000101111010010000011110;
         rom[1358] = 24'b000101111111100001101001;
         rom[1359] = 24'b000110000011000101010110;
         rom[1360] = 24'b000110001011011010101010;
         rom[1361] = 24'b000110100100101001001011;
         rom[1362] = 24'b000110101111000101001011;
         rom[1363] = 24'b000110110110111011010100;
         rom[1364] = 24'b000111000001011111111000;
         rom[1365] = 24'b000111001010010111011111;
         rom[1366] = 24'b000111010011111110011111;
         rom[1367] = 24'b000111100010111010110100;
         rom[1368] = 24'b001000001000101100100010;
         rom[1369] = 24'b001000000101101110111100;
         rom[1370] = 24'b001000010111110100110110;
         rom[1371] = 24'b001000011110100001110101;
         rom[1372] = 24'b001000100111111100100000;
         rom[1373] = 24'b001001000000001001000111;
         rom[1374] = 24'b001000111011101001000010;
         rom[1375] = 24'b001001010110110101010100;
         rom[1376] = 24'b001001001001000111001000;
         rom[1377] = 24'b001001000100110110001100;
         rom[1378] = 24'b001001010010111000111010;
         rom[1379] = 24'b001001010011011011000101;
         rom[1380] = 24'b001001100011100001110101;
         rom[1381] = 24'b001001100000011110100001;
         rom[1382] = 24'b001001011001000000000100;
         rom[1383] = 24'b001001011111010100110010;
         rom[1384] = 24'b001001100001101111100100;
         rom[1385] = 24'b001001011110001101001111;
         rom[1386] = 24'b001001100110011000100011;
         rom[1387] = 24'b001001100101010001011011;
         rom[1388] = 24'b001001100001010111100010;
         rom[1389] = 24'b001001010000100101101111;
         rom[1390] = 24'b001001001110011000101100;
         rom[1391] = 24'b001000110101111111100011;
         rom[1392] = 24'b001000110111001011001010;
         rom[1393] = 24'b001000101010101101010001;
         rom[1394] = 24'b001000101001100101011010;
         rom[1395] = 24'b001000110001100101001000;
         rom[1396] = 24'b001000101000100111011110;
         rom[1397] = 24'b001000101100101000001010;
         rom[1398] = 24'b001000100110100001101011;
         rom[1399] = 24'b001000011101111111110111;
         rom[1400] = 24'b001000100010100001010011;
         rom[1401] = 24'b001000010111011100100001;
         rom[1402] = 24'b001000010101100001110101;
         rom[1403] = 24'b001000110010000111001010;
         rom[1404] = 24'b001000011001010100010001;
         rom[1405] = 24'b001000011110000111100100;
         rom[1406] = 24'b001000001111011010111001;
         rom[1407] = 24'b001000011010001101101101;
         rom[1408] = 24'b001000010010000000100101;
         rom[1409] = 24'b001000001100010001001110;
         rom[1410] = 24'b000111111110010100100010;
         rom[1411] = 24'b000111101011001001000111;
         rom[1412] = 24'b000111110111111101110111;
         rom[1413] = 24'b000111001110100010010110;
         rom[1414] = 24'b000111001001010101011001;
         rom[1415] = 24'b000111000111110111011010;
         rom[1416] = 24'b000110110001111010011011;
         rom[1417] = 24'b000110101011001101101010;
         rom[1418] = 24'b000110011100111001101011;
         rom[1419] = 24'b000110000011110101111110;
         rom[1420] = 24'b000110000011010100000110;
         rom[1421] = 24'b000101101101111111011110;
         rom[1422] = 24'b000101011100101011111100;
         rom[1423] = 24'b000101100001000101111111;
         rom[1424] = 24'b000101011001000011110101;
         rom[1425] = 24'b000101001101011111001100;
         rom[1426] = 24'b000101000010000100001110;
         rom[1427] = 24'b000100110011101100001110;
         rom[1428] = 24'b000100111100110110000011;
         rom[1429] = 24'b000100111000111011111010;
         rom[1430] = 24'b000100110001110011001110;
         rom[1431] = 24'b000100110000110100011100;
         rom[1432] = 24'b000100110101001000011111;
         rom[1433] = 24'b000100101110001010100110;
         rom[1434] = 24'b000100110011101110111001;
         rom[1435] = 24'b000100110000011100111010;
         rom[1436] = 24'b000100110001110001100110;
         rom[1437] = 24'b000100101110110000100110;
         rom[1438] = 24'b000100101101111110001000;
         rom[1439] = 24'b000100101010010000011011;
         rom[1440] = 24'b000100101011101111101000;
         rom[1441] = 24'b000100101000110110111100;
         rom[1442] = 24'b000100011101100110010101;
         rom[1443] = 24'b000100001001000011100101;
         rom[1444] = 24'b000100000010010010111101;
         rom[1445] = 24'b000011110011100001100111;
         rom[1446] = 24'b000011110011010001010000;
         rom[1447] = 24'b000011100001010000010010;
         rom[1448] = 24'b000011011100000111111110;
         rom[1449] = 24'b000010111110101010110101;
         rom[1450] = 24'b000010111101011101101111;
         rom[1451] = 24'b000010101101001000001010;
         rom[1452] = 24'b000010001110010011010000;
         rom[1453] = 24'b000010011100001100010100;
         rom[1454] = 24'b000010000101001110010100;
         rom[1455] = 24'b000001111001001011010100;
         rom[1456] = 24'b000001101010101011000101;
         rom[1457] = 24'b000001100010100010000011;
         rom[1458] = 24'b000001011001011111111000;
         rom[1459] = 24'b000001001000111011101100;
         rom[1460] = 24'b000001000010111011100010;
         rom[1461] = 24'b000001000010101000000010;
         rom[1462] = 24'b000001010101101011001110;
         rom[1463] = 24'b000001000110011011110010;
         rom[1464] = 24'b000001000101101110001000;
         rom[1465] = 24'b000000111101100000010101;
         rom[1466] = 24'b000001000101101101101010;
         rom[1467] = 24'b000001000010100011110000;
         rom[1468] = 24'b000000110101110110101101;
         rom[1469] = 24'b000001000001000111110001;
         rom[1470] = 24'b000001000000111100101100;
         rom[1471] = 24'b000000101110010110010000;
         rom[1472] = 24'b000000111001000101011111;
         rom[1473] = 24'b000000100101001101001011;
         rom[1474] = 24'b000000101000101010111000;
         rom[1475] = 24'b000000011110111010011110;
         rom[1476] = 24'b000000011110010111100110;
         rom[1477] = 24'b000000011100101101111000;
         rom[1478] = 24'b000000010000100100001001;
         rom[1479] = 24'b000000000110001011110100;
         rom[1480] = 24'b111111101110110010100011;
         rom[1481] = 24'b111111011111100010101110;
         rom[1482] = 24'b111111100001111110111010;
         rom[1483] = 24'b111111001101010000110100;
         rom[1484] = 24'b111110111011011111100010;
         rom[1485] = 24'b111110110001010000000000;
         rom[1486] = 24'b111110010000100001000011;
         rom[1487] = 24'b111110010010101110000100;
         rom[1488] = 24'b111110001110010100001001;
         rom[1489] = 24'b111110010101001010110111;
         rom[1490] = 24'b111110001110101010011111;
         rom[1491] = 24'b111110010110111010011010;
         rom[1492] = 24'b111110101001001100110111;
         rom[1493] = 24'b111110101010110110011010;
         rom[1494] = 24'b111110101111010101001001;
         rom[1495] = 24'b111111000001111101110000;
         rom[1496] = 24'b111110111100011111000110;
         rom[1497] = 24'b111111010101010001010100;
         rom[1498] = 24'b111111100011011100111100;
         rom[1499] = 24'b111111101111101000111110;
         rom[1500] = 24'b111111111110000101001010;
         rom[1501] = 24'b000000000100111001010100;
         rom[1502] = 24'b000000010100010001101110;
         rom[1503] = 24'b000000010111101001111110;
         rom[1504] = 24'b000000011110011100111001;
         rom[1505] = 24'b000000100000100000101101;
         rom[1506] = 24'b000000011000111010110011;
         rom[1507] = 24'b000000101111010111011101;
         rom[1508] = 24'b000000010100111110011000;
         rom[1509] = 24'b000000101010111110101010;
         rom[1510] = 24'b000000100100110100110001;
         rom[1511] = 24'b000000011001001100010011;
         rom[1512] = 24'b000000011101111001111010;
         rom[1513] = 24'b000000011110010010010011;
         rom[1514] = 24'b000000001011110111100110;
         rom[1515] = 24'b000000001111011001101000;
         rom[1516] = 24'b000000000010101100001001;
         rom[1517] = 24'b111111111000001010000101;
         rom[1518] = 24'b111111111011000101010110;
         rom[1519] = 24'b111111110011101001101111;
         rom[1520] = 24'b111111101011010111111110;
         rom[1521] = 24'b111111101011111111001011;
         rom[1522] = 24'b111111101001010011101001;
         rom[1523] = 24'b111111011101011010000011;
         rom[1524] = 24'b111111010111010010000110;
         rom[1525] = 24'b111111011110001100010110;
         rom[1526] = 24'b111111011000110110011111;
         rom[1527] = 24'b111111011000100110001000;
         rom[1528] = 24'b111111100010011111110100;
         rom[1529] = 24'b111111011101100110101011;
         rom[1530] = 24'b111111111001000100100111;
         rom[1531] = 24'b111111111010000000101111;
         rom[1532] = 24'b111111111000010011110100;
         rom[1533] = 24'b111111111101111010100000;
         rom[1534] = 24'b000000000011000110000100;
         rom[1535] = 24'b000000010011100100011010;
         rom[1536] = 24'b000000010010011010100000;
         rom[1537] = 24'b000000010010001010011111;
         rom[1538] = 24'b000000011001100000101110;
         rom[1539] = 24'b000000100101001100100110;
         rom[1540] = 24'b000000101010100010101000;
         rom[1541] = 24'b000000100011011000110011;
         rom[1542] = 24'b000000100001101101100110;
         rom[1543] = 24'b000000100001101010110110;
         rom[1544] = 24'b000000101010010001010011;
         rom[1545] = 24'b000000001111101100101010;
         rom[1546] = 24'b000000011001001001011100;
         rom[1547] = 24'b000000011001011010100110;
         rom[1548] = 24'b111111111110001111111100;
         rom[1549] = 24'b000000001010100000000100;
         rom[1550] = 24'b000000000110001000010000;
         rom[1551] = 24'b111111100111110011001000;
         rom[1552] = 24'b111111101101010001010001;
         rom[1553] = 24'b111111100111000010101100;
         rom[1554] = 24'b111111011010101110100010;
         rom[1555] = 24'b111111100010010111011111;
         rom[1556] = 24'b111111100011101001010010;
         rom[1557] = 24'b111111100101111101011111;
         rom[1558] = 24'b111111101101111100100001;
         rom[1559] = 24'b111111101000100111111101;
         rom[1560] = 24'b111111011000001000001111;
         rom[1561] = 24'b111111011010110110010010;
         rom[1562] = 24'b111111100111100100011110;
         rom[1563] = 24'b111111101001001011001111;
         rom[1564] = 24'b111111110100110001010111;
         rom[1565] = 24'b111111110010011010100001;
         rom[1566] = 24'b111111110110111000011100;
         rom[1567] = 24'b000000000100101001001110;
         rom[1568] = 24'b111111111101011010001010;
         rom[1569] = 24'b000000001111010010000100;
         rom[1570] = 24'b000000011011101110100110;
         rom[1571] = 24'b000000100010011011101010;
         rom[1572] = 24'b000000011010100110001010;
         rom[1573] = 24'b000000100101010100100111;
         rom[1574] = 24'b000000100111011110110111;
         rom[1575] = 24'b000000100100111110010011;
         rom[1576] = 24'b000000011101001001101100;
         rom[1577] = 24'b000000010111111001111111;
         rom[1578] = 24'b000000010101100011001101;
         rom[1579] = 24'b000000011110001110100001;
         rom[1580] = 24'b000000011101111000001000;
         rom[1581] = 24'b000000010101100111111111;
         rom[1582] = 24'b000000001011110101010000;
         rom[1583] = 24'b111111111010011011110111;
         rom[1584] = 24'b111111111000100001110111;
         rom[1585] = 24'b111111110011111101010001;
         rom[1586] = 24'b111111100100111010000001;
         rom[1587] = 24'b111111101011000111110111;
         rom[1588] = 24'b111111101011101011110010;
         rom[1589] = 24'b111111010100101010100101;
         rom[1590] = 24'b111111011100010110011110;
         rom[1591] = 24'b111111011111011001010011;
         rom[1592] = 24'b111111010111111110000111;
         rom[1593] = 24'b111111011010110011000100;
         rom[1594] = 24'b111111101001101111100100;
         rom[1595] = 24'b111111100001001111010111;
         rom[1596] = 24'b111111100110111110100110;
         rom[1597] = 24'b000000000001000001000110;
         rom[1598] = 24'b111111101000011101111000;
         rom[1599] = 24'b111111110011101100000101;
         rom[1600] = 24'b111111110110111000011101;
         rom[1601] = 24'b000000000100111010011010;
         rom[1602] = 24'b000000010111000101011100;
         rom[1603] = 24'b000000010010000101000001;
         rom[1604] = 24'b000000011000100101110100;
         rom[1605] = 24'b000000100010000110010110;
         rom[1606] = 24'b000000011111011011010000;
         rom[1607] = 24'b000000101011101011001010;
         rom[1608] = 24'b000000100111000101101010;
         rom[1609] = 24'b000000100010100011010010;
         rom[1610] = 24'b000000011010110101001001;
         rom[1611] = 24'b000000011101000011110100;
         rom[1612] = 24'b000000010010000101111001;
         rom[1613] = 24'b000000010000001110010000;
         rom[1614] = 24'b000000000110001101110101;
         rom[1615] = 24'b000000001001111101010100;
         rom[1616] = 24'b000000000011100111100000;
         rom[1617] = 24'b111111111001000111001111;
         rom[1618] = 24'b111111110001011111110101;
         rom[1619] = 24'b111111110101011100110001;
         rom[1620] = 24'b111111101001000010001101;
         rom[1621] = 24'b111111101111101010000011;
         rom[1622] = 24'b111111100010001000100111;
         rom[1623] = 24'b111111101010111001110110;
         rom[1624] = 24'b111111100000000110100011;
         rom[1625] = 24'b111111100000000100100111;
         rom[1626] = 24'b111111011110111111001101;
         rom[1627] = 24'b111111101010110110010010;
         rom[1628] = 24'b111111101101101010101111;
         rom[1629] = 24'b111111100111001101001001;
         rom[1630] = 24'b111111101001100000001100;
         rom[1631] = 24'b111111101101000110101101;
         rom[1632] = 24'b000000000010011000110101;
         rom[1633] = 24'b000000001010110000100110;
         rom[1634] = 24'b111111111111101000000010;
         rom[1635] = 24'b111111111000111101111001;
         rom[1636] = 24'b000000001001010001111111;
         rom[1637] = 24'b000000100011010000110110;
         rom[1638] = 24'b000000011000011001111101;
         rom[1639] = 24'b000000100001111000101000;
         rom[1640] = 24'b000000100001000000010000;
         rom[1641] = 24'b000000101111111001110010;
         rom[1642] = 24'b000000110110000101111001;
         rom[1643] = 24'b000000101001111101000101;
         rom[1644] = 24'b000000111000100111111110;
         rom[1645] = 24'b000001000010001011110001;
         rom[1646] = 24'b000000110111111100011000;
         rom[1647] = 24'b000000110011110011001011;
         rom[1648] = 24'b000000011110100110010001;
         rom[1649] = 24'b000000101100000100101011;
         rom[1650] = 24'b000000101010011010110111;
         rom[1651] = 24'b000000101001101110010000;
         rom[1652] = 24'b000000100010001100101111;
         rom[1653] = 24'b000000010111101100001000;
         rom[1654] = 24'b000000011100000100000111;
         rom[1655] = 24'b000000001110101100100100;
         rom[1656] = 24'b000000010010101011000110;
         rom[1657] = 24'b000000001000001111000000;
         rom[1658] = 24'b000000001001000011000011;
         rom[1659] = 24'b000000010110010011001000;
         rom[1660] = 24'b000000001101110111001011;
         rom[1661] = 24'b000000011101000101111011;
         rom[1662] = 24'b000000010101100110011011;
         rom[1663] = 24'b000000011111010001111101;
         rom[1664] = 24'b000000101101010101011001;
         rom[1665] = 24'b000000100010000110100111;
         rom[1666] = 24'b000000110101001000000000;
         rom[1667] = 24'b000001001101100100110010;
         rom[1668] = 24'b000001000000010110010101;
         rom[1669] = 24'b000001100100110010001011;
         rom[1670] = 24'b000001010110000001101001;
         rom[1671] = 24'b000001011011111110111001;
         rom[1672] = 24'b000001011110000011001010;
         rom[1673] = 24'b000001100000000010000110;
         rom[1674] = 24'b000001101010110011100111;
         rom[1675] = 24'b000001101100000001101011;
         rom[1676] = 24'b000001110100000010110010;
         rom[1677] = 24'b000001101001001010111100;
         rom[1678] = 24'b000001101001001101011000;
         rom[1679] = 24'b000001011100111110101011;
         rom[1680] = 24'b000001100010101000110111;
         rom[1681] = 24'b000001101001010101111101;
         rom[1682] = 24'b000001010010111100110000;
         rom[1683] = 24'b000001000000011110000110;
         rom[1684] = 24'b000001000110111011111001;
         rom[1685] = 24'b000000110010100001101010;
         rom[1686] = 24'b000000110100101010010100;
         rom[1687] = 24'b000001000001110001100010;
         rom[1688] = 24'b000000101011101001011111;
         rom[1689] = 24'b000000110110011000001100;
         rom[1690] = 24'b000000110101100001011011;
         rom[1691] = 24'b000000110111101011000101;
         rom[1692] = 24'b000000110011010000011101;
         rom[1693] = 24'b000000101011001001111101;
         rom[1694] = 24'b000000111010011011001011;
         rom[1695] = 24'b000000111101100100011001;
         rom[1696] = 24'b000001000001110111101010;
         rom[1697] = 24'b000001000111111011001100;
         rom[1698] = 24'b000001001000110111010111;
         rom[1699] = 24'b000001011001100110100011;
         rom[1700] = 24'b000001011001110010000111;
         rom[1701] = 24'b000001101101100000100001;
         rom[1702] = 24'b000001101010111011111010;
         rom[1703] = 24'b000001101110100111011110;
         rom[1704] = 24'b000001111110000000001000;
         rom[1705] = 24'b000001110100101001101000;
         rom[1706] = 24'b000010000001101101110011;
         rom[1707] = 24'b000010000100000010100001;
         rom[1708] = 24'b000010000000110001000110;
         rom[1709] = 24'b000010010000010000111001;
         rom[1710] = 24'b000010001011111000101001;
         rom[1711] = 24'b000010001010011110110001;
         rom[1712] = 24'b000001110110101101101010;
         rom[1713] = 24'b000001111111111111110011;
         rom[1714] = 24'b000001111011001100010011;
         rom[1715] = 24'b000001111111101111001111;
         rom[1716] = 24'b000001101010111101010001;
         rom[1717] = 24'b000001011100101010101111;
         rom[1718] = 24'b000001010100011101100101;
         rom[1719] = 24'b000001010011011000011011;
         rom[1720] = 24'b000001001111001100000000;
         rom[1721] = 24'b000001001100100000000101;
         rom[1722] = 24'b000001001011000000101111;
         rom[1723] = 24'b000001000001001110011101;
         rom[1724] = 24'b000000111110111101100111;
         rom[1725] = 24'b000001000001100010101111;
         rom[1726] = 24'b000000111011000001010111;
         rom[1727] = 24'b000000111100101000101010;
         rom[1728] = 24'b000001010100000011010010;
         rom[1729] = 24'b000001001110101011110100;
         rom[1730] = 24'b000001011101110110011010;
         rom[1731] = 24'b000001011000110001110011;
         rom[1732] = 24'b000001100010101101100011;
         rom[1733] = 24'b000001101001111111100000;
         rom[1734] = 24'b000001101010111001000011;
         rom[1735] = 24'b000010000100010111010010;
         rom[1736] = 24'b000001111010101011100101;
         rom[1737] = 24'b000001111101000101101000;
         rom[1738] = 24'b000010000010100000001000;
         rom[1739] = 24'b000010000111001111010011;
         rom[1740] = 24'b000010001000001010100000;
         rom[1741] = 24'b000010011001101000111001;
         rom[1742] = 24'b000010010001101000010101;
         rom[1743] = 24'b000010100011110101000101;
         rom[1744] = 24'b000010001110101100101110;
         rom[1745] = 24'b000010011000101100101101;
         rom[1746] = 24'b000010000010110100001010;
         rom[1747] = 24'b000010000101011001000101;
         rom[1748] = 24'b000001110111101001110111;
         rom[1749] = 24'b000001110001011011001010;
         rom[1750] = 24'b000001101010111011000101;
         rom[1751] = 24'b000001101001100011000001;
         rom[1752] = 24'b000001101001001001111010;
         rom[1753] = 24'b000001011011010000110100;
         rom[1754] = 24'b000001001000100110100110;
         rom[1755] = 24'b000001000111001011101001;
         rom[1756] = 24'b000001010000010011010110;
         rom[1757] = 24'b000001000010101101010110;
         rom[1758] = 24'b000001010101100101010001;
         rom[1759] = 24'b000001011101110010101010;
         rom[1760] = 24'b000001001001000110010010;
         rom[1761] = 24'b000001100000111101101001;
         rom[1762] = 24'b000001011000110011110110;
         rom[1763] = 24'b000001010011110010101110;
         rom[1764] = 24'b000001010110111110010011;
         rom[1765] = 24'b000001101011011010111000;
         rom[1766] = 24'b000001100110000000101100;
         rom[1767] = 24'b000001110010010111011011;
         rom[1768] = 24'b000010000000111011011001;
         rom[1769] = 24'b000010000101010011101010;
         rom[1770] = 24'b000010001011000010000110;
         rom[1771] = 24'b000010011000100011000110;
         rom[1772] = 24'b000010011010111100001100;
         rom[1773] = 24'b000010001101101010000001;
         rom[1774] = 24'b000010100011110110111101;
         rom[1775] = 24'b000010011100100011000011;
         rom[1776] = 24'b000010011011110101001001;
         rom[1777] = 24'b000010011110110011100001;
         rom[1778] = 24'b000010010000100001111111;
         rom[1779] = 24'b000010001011111011101100;
         rom[1780] = 24'b000010011011100100100001;
         rom[1781] = 24'b000010001010000110110100;
         rom[1782] = 24'b000001111011011110110000;
         rom[1783] = 24'b000001110000010001010101;
         rom[1784] = 24'b000010000011111001111101;
         rom[1785] = 24'b000001101010011001011001;
         rom[1786] = 24'b000001100100011001111001;
         rom[1787] = 24'b000001010100010011010111;
         rom[1788] = 24'b000001010101001101100100;
         rom[1789] = 24'b000001010100001011111011;
         rom[1790] = 24'b000001100001011001010011;
         rom[1791] = 24'b000001010000101011010001;
         rom[1792] = 24'b000001010101001010101111;
         rom[1793] = 24'b000001010100001100000001;
         rom[1794] = 24'b000001010001100011000000;
         rom[1795] = 24'b000001011010010001101001;
         rom[1796] = 24'b000001011010100000110000;
         rom[1797] = 24'b000001101011011100011010;
         rom[1798] = 24'b000001100010111000000100;
         rom[1799] = 24'b000001101010010010000001;
         rom[1800] = 24'b000001110101001001110111;
         rom[1801] = 24'b000001111101101011011000;
         rom[1802] = 24'b000010000001000010111110;
         rom[1803] = 24'b000010001101000111010100;
         rom[1804] = 24'b000010010010101010010101;
         rom[1805] = 24'b000010010001011010010111;
         rom[1806] = 24'b000010010010100011111110;
         rom[1807] = 24'b000010101010110100010001;
         rom[1808] = 24'b000010100111110011100100;
         rom[1809] = 24'b000010100000010011010000;
         rom[1810] = 24'b000010010100100101101100;
         rom[1811] = 24'b000010011011000000110100;
         rom[1812] = 24'b000010100010010100110111;
         rom[1813] = 24'b000010000101000011100101;
         rom[1814] = 24'b000010000011100110101110;
         rom[1815] = 24'b000010000010010101001010;
         rom[1816] = 24'b000010000100010111110000;
         rom[1817] = 24'b000001110111001111010111;
         rom[1818] = 24'b000001100100101000001100;
         rom[1819] = 24'b000001110010110111100011;
         rom[1820] = 24'b000001010000010100110001;
         rom[1821] = 24'b000001100110011011111000;
         rom[1822] = 24'b000001100110001010110101;
         rom[1823] = 24'b000001011101011001000110;
         rom[1824] = 24'b000001001111100100100111;
         rom[1825] = 24'b000001011000110001110110;
         rom[1826] = 24'b000001011100110010001110;
         rom[1827] = 24'b000001001010010011111101;
         rom[1828] = 24'b000001001001101110110110;
         rom[1829] = 24'b000001100111111101111001;
         rom[1830] = 24'b000001011001100010000111;
         rom[1831] = 24'b000001101010110011000100;
         rom[1832] = 24'b000001101100001100010111;
         rom[1833] = 24'b000001110111010100000010;
         rom[1834] = 24'b000001110011100010110000;
         rom[1835] = 24'b000010000001011001000001;
         rom[1836] = 24'b000010001011100000001101;
         rom[1837] = 24'b000010001111011010000111;
         rom[1838] = 24'b000010011011111011000111;
         rom[1839] = 24'b000010100110101101100111;
         rom[1840] = 24'b000010011000110000101110;
         rom[1841] = 24'b000010011111010010100010;
         rom[1842] = 24'b000010011101001011100000;
         rom[1843] = 24'b000010011010000100111100;
         rom[1844] = 24'b000010011110000110010110;
         rom[1845] = 24'b000010001100001011001001;
         rom[1846] = 24'b000010011101110100100110;
         rom[1847] = 24'b000010001110111100111000;
         rom[1848] = 24'b000001110111100001111111;
         rom[1849] = 24'b000001111101110110001001;
         rom[1850] = 24'b000001111011000010111000;
         rom[1851] = 24'b000001101001010101010011;
         rom[1852] = 24'b000001111010100001100010;
         rom[1853] = 24'b000001011110010001110100;
         rom[1854] = 24'b000001010100100010101011;
         rom[1855] = 24'b000001011110010001101111;
         rom[1856] = 24'b000001010000111100011101;
         rom[1857] = 24'b000001010100011001000000;
         rom[1858] = 24'b000001010100000100001001;
         rom[1859] = 24'b000001011001010111111100;
         rom[1860] = 24'b000001010001010011111000;
         rom[1861] = 24'b000001011100101100011001;
         rom[1862] = 24'b000001010100100100111111;
         rom[1863] = 24'b000001011000010011101010;
         rom[1864] = 24'b000001101001000000111000;
         rom[1865] = 24'b000001101010101001000101;
         rom[1866] = 24'b000001101001011011001101;
         rom[1867] = 24'b000001111100101101000110;
         rom[1868] = 24'b000010001000011001100001;
         rom[1869] = 24'b000010000111001110110011;
         rom[1870] = 24'b000010001101001111101110;
         rom[1871] = 24'b000010000101000100001100;
         rom[1872] = 24'b000010011010101101101001;
         rom[1873] = 24'b000010011010001010001011;
         rom[1874] = 24'b000010011111001001111101;
         rom[1875] = 24'b000010001100101100110101;
         rom[1876] = 24'b000010100101000001110001;
         rom[1877] = 24'b000010100110101011001010;
         rom[1878] = 24'b000010010101100110011000;
         rom[1879] = 24'b000010011110111110111000;
         rom[1880] = 24'b000010010000101101110101;
         rom[1881] = 24'b000010000111111101110100;
         rom[1882] = 24'b000001110110101001101110;
         rom[1883] = 24'b000001111010001110110000;
         rom[1884] = 24'b000001111001110001011101;
         rom[1885] = 24'b000001100010001000010010;
         rom[1886] = 24'b000001011110011010111110;
         rom[1887] = 24'b000001100011111110000001;
         rom[1888] = 24'b000001011000101111000010;
         rom[1889] = 24'b000001001001110010101100;
         rom[1890] = 24'b000001011100111100010111;
         rom[1891] = 24'b000001000100011101001101;
         rom[1892] = 24'b000001001101100100000000;
         rom[1893] = 24'b000001000001010011111101;
         rom[1894] = 24'b000001010100010100001010;
         rom[1895] = 24'b000001011000101101111110;
         rom[1896] = 24'b000001001100000110011100;
         rom[1897] = 24'b000001001100111100011000;
         rom[1898] = 24'b000001011001101010000010;
         rom[1899] = 24'b000001100111011110011011;
         rom[1900] = 24'b000001101010000001011000;
         rom[1901] = 24'b000001101110010010001011;
         rom[1902] = 24'b000010000001001101111110;
         rom[1903] = 24'b000010000101010101101110;
         rom[1904] = 24'b000001110100010000010011;
         rom[1905] = 24'b000010010001100011110101;
         rom[1906] = 24'b000010001111110100010110;
         rom[1907] = 24'b000010011011010011010111;
         rom[1908] = 24'b000010000101101001011000;
         rom[1909] = 24'b000010001011101000011100;
         rom[1910] = 24'b000010000110011011110000;
         rom[1911] = 24'b000010001101011010101000;
         rom[1912] = 24'b000001111101001110100110;
         rom[1913] = 24'b000010000110001101010100;
         rom[1914] = 24'b000001110011100110011110;
         rom[1915] = 24'b000001110110001111110100;
         rom[1916] = 24'b000001101000010111111111;
         rom[1917] = 24'b000001011101101000111100;
         rom[1918] = 24'b000001001110011111000101;
         rom[1919] = 24'b000001010011001110110011;
         rom[1920] = 24'b000001001101110100100001;
         rom[1921] = 24'b000001001101011101000001;
         rom[1922] = 24'b000000111000011100000010;
         rom[1923] = 24'b000001000110110010011000;
         rom[1924] = 24'b000001001000101101010011;
         rom[1925] = 24'b000001000110011011101011;
         rom[1926] = 24'b000001000100001000011101;
         rom[1927] = 24'b000000111101111111100011;
         rom[1928] = 24'b000000110001010101011100;
         rom[1929] = 24'b000001000111010000001101;
         rom[1930] = 24'b000001010001111011001110;
         rom[1931] = 24'b000001010011001101110111;
         rom[1932] = 24'b000001010111110101001101;
         rom[1933] = 24'b000001010100011000101000;
         rom[1934] = 24'b000001101010111111111100;
         rom[1935] = 24'b000001110101100110111110;
         rom[1936] = 24'b000001111011000001010100;
         rom[1937] = 24'b000001110000100111101100;
         rom[1938] = 24'b000010000001011010101001;
         rom[1939] = 24'b000001111000011001011100;
         rom[1940] = 24'b000001111011110010010100;
         rom[1941] = 24'b000001111011100111111000;
         rom[1942] = 24'b000001111000100101101011;
         rom[1943] = 24'b000010000010100101010111;
         rom[1944] = 24'b000010000111010000100000;
         rom[1945] = 24'b000001101101110011001100;
         rom[1946] = 24'b000001100101000110011000;
         rom[1947] = 24'b000001101000111001110111;
         rom[1948] = 24'b000001100110100101010001;
         rom[1949] = 24'b000001011001000110010011;
         rom[1950] = 24'b000001010010111100110011;
         rom[1951] = 24'b000001011101100000110100;
         rom[1952] = 24'b000001000011100101001010;
         rom[1953] = 24'b000000111010101010101001;
         rom[1954] = 24'b000000110111111001110010;
         rom[1955] = 24'b000000110001000001100111;
         rom[1956] = 24'b000000100010000101101111;
         rom[1957] = 24'b000000101111111110111001;
         rom[1958] = 24'b000000101101110110100011;
         rom[1959] = 24'b000000111000010100001101;
         rom[1960] = 24'b000000100010110000010010;
         rom[1961] = 24'b000000101101001111111110;
         rom[1962] = 24'b000000101100001000011000;
         rom[1963] = 24'b000000110111110100110100;
         rom[1964] = 24'b000000111011101100001011;
         rom[1965] = 24'b000000100111100011111010;
         rom[1966] = 24'b000000111010010110001100;
         rom[1967] = 24'b000001001011001010011000;
         rom[1968] = 24'b000001001110011010100111;
         rom[1969] = 24'b000001010100101110001110;
         rom[1970] = 24'b000001011101010110100111;
         rom[1971] = 24'b000001100110011010010011;
         rom[1972] = 24'b000001010100100101111001;
         rom[1973] = 24'b000001100010110111011101;
         rom[1974] = 24'b000001101010011110111001;
         rom[1975] = 24'b000001101100010100010101;
         rom[1976] = 24'b000001101001011010000100;
         rom[1977] = 24'b000001100110110010001100;
         rom[1978] = 24'b000001010011100010001110;
         rom[1979] = 24'b000001001110111011101011;
         rom[1980] = 24'b000001001011100010000110;
         rom[1981] = 24'b000001000100101011100010;
         rom[1982] = 24'b000000111001110000001110;
         rom[1983] = 24'b000000110011101000100011;
         rom[1984] = 24'b000000101111000110011010;
         rom[1985] = 24'b000000101001111111111110;
         rom[1986] = 24'b000000100111101100011011;
         rom[1987] = 24'b000000010100110101001101;
         rom[1988] = 24'b111111111111101101101010;
         rom[1989] = 24'b111111111111101000110111;
         rom[1990] = 24'b111111110110000111000100;
         rom[1991] = 24'b000000001100011100111101;
         rom[1992] = 24'b111111110101101010010001;
         rom[1993] = 24'b000000001011111010101001;
         rom[1994] = 24'b111111110100100110110011;
         rom[1995] = 24'b000000000110100111110111;
         rom[1996] = 24'b111111111010011011011010;
         rom[1997] = 24'b000000001111001001000101;
         rom[1998] = 24'b111111111110111010011100;
         rom[1999] = 24'b000000000001010001110000;
         end 

	 always @(posedge(clk))
		 begin 
			 if(reset) 
				 begin 
					 data_out <= 24'b0; 
					 i <= 16'b0; 
					 counter <= 16'b0; 
				 end 
			 else 
				 begin 
					 if(counter == 16'd5000) 
						 begin 
							 data_out <= rom[i]; 
							 counter <=16'b0; 
							 if(i == 1999) i <= 0; 
							 else i <= i + 1; 
						 end 
					 else counter <= counter + 16'd1; 
				 end 
		 end 

endmodule
