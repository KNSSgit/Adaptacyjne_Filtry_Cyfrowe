//////////////////////////////////////////////////////////////////////////////////
// Kolo Naukowe Systemow Scalonych
// 10.2017
// 
// Modul: gen_sinus_zabrudzony
// Projekt: Adaptacyjne filtry cyfrowe do kondycjonowania sygnalow biomedycznych 
// Model urzadzenia: Nexys Video Artix 7 (XC7A200T-1SBG484C)
// 
// Wersja: 0.1
//////////////////////////////////////////////////////////////////////////////////


module gen_sinus_zabrudzony(
    output reg signed [23:0] data_out,
    input clk,
    input reset
    );
    
    reg signed [23:0] rom [0:39];
    reg [8:0] i;
    reg [15:0] counter;//50000 * 40pr�bek = 2 000 000 ; zegar 100mhz => 50hz

    always @(reset)
        begin
        rom[0] = 24'b000000000000000000000000;
        rom[1] = 24'b001001100111101011101000;
        rom[2] = 24'b010000110000100111101101;
        rom[3] = 24'b010011110110110100111001;
        rom[4] = 24'b010010110101011010110100;
        rom[5] = 24'b001111000110101111110110;
        rom[6] = 24'b001011000000010001011000;
        rom[7] = 24'b001000111000000010010110;
        rom[8] = 24'b001010001010001000101110;
        rom[9] = 24'b001110110100100011001000;
        rom[10] = 24'b010101010111001100000000;
        rom[11] = 24'b011011011000001010010101;
        rom[12] = 24'b011110011110011010001011;
        rom[13] = 24'b011101001100010011110011;
        rom[14] = 24'b010111100011111000100110;
        rom[15] = 24'b001111000110101111110110;
        rom[16] = 24'b000110010001110011100111;
        rom[17] = 24'b111111100010100011011101;
        rom[18] = 24'b111100011100010110010001;
        rom[19] = 24'b111101000100000100011010;
        rom[20] = 24'b000000000000000000000000;
        rom[21] = 24'b000010111011111011100110;
        rom[22] = 24'b000011100011101001101111;
        rom[23] = 24'b000000011101011100100011;
        rom[24] = 24'b111001101110001100011001;
        rom[25] = 24'b110000111001010000001010;
        rom[26] = 24'b101000011100000111011010;
        rom[27] = 24'b100010110011101100001101;
        rom[28] = 24'b100001100001100101110101;
        rom[29] = 24'b100100100111110101101011;
        rom[30] = 24'b101010101000110100000000;
        rom[31] = 24'b110001001011011100111000;
        rom[32] = 24'b110101110101110111010010;
        rom[33] = 24'b110111000111111101101010;
        rom[34] = 24'b110100111111101110101000;
        rom[35] = 24'b110000111001010000001010;
        rom[36] = 24'b101101001010100101001100;
        rom[37] = 24'b101100001001001011000111;
        rom[38] = 24'b101111001111011000010011;
        rom[39] = 24'b110110011000010100011000;

        end
        
        always @(posedge(clk))
            begin
                if(reset)
                    begin
                        data_out <= 24'b0;
                        i <= 9'b0;
                        counter <= 16'b0;
                    end
                else
                    begin
                        if(counter == 16'd50000)
                            begin
                                data_out <= rom[i];
                                counter <= 16'b0;
                                if(i == 39) i <= 0;
                                else i <= i + 1;
                            end
                        else counter <= counter + 16'd1;
                    end
            end
            
endmodule
