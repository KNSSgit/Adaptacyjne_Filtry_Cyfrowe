module gen_ekg_55(
 	 output reg signed [23:0] data_out,
	 input clk,
	 input reset
	 ); 

	 reg signed [23:0] rom[0:1999];
	 reg [15:0] i;
	 reg [15:0] counter;//5000 * 2000pr�bek = 10 000 000 ; zegar 10mhz => 1hz

	 always @(reset)     // fs = 2kHz; f1 = 1Hz; A1 = 3000000; f2 = 55Hz; A2 = 150000
		 begin 
         rom[0] = 24'b111111110101110110001110;
         rom[1] = 24'b000000000011110000011111;
         rom[2] = 24'b000000001110010010011010;
         rom[3] = 24'b000000001110111110010100;
         rom[4] = 24'b000000011000001001101000;
         rom[5] = 24'b000000010000111111010100;
         rom[6] = 24'b000000010100101001110000;
         rom[7] = 24'b000000100111010110101111;
         rom[8] = 24'b000000011110101101010100;
         rom[9] = 24'b000000011011000110101001;
         rom[10] = 24'b000000101011101110111001;
         rom[11] = 24'b000000101010100011010000;
         rom[12] = 24'b000000011101000000101001;
         rom[13] = 24'b000000011101010111000001;
         rom[14] = 24'b000000101011001001001110;
         rom[15] = 24'b000000001101100101101000;
         rom[16] = 24'b000000001100111010101100;
         rom[17] = 24'b000000001000001111011111;
         rom[18] = 24'b111111111101000011010101;
         rom[19] = 24'b111111111101011111001100;
         rom[20] = 24'b111111101100110001011101;
         rom[21] = 24'b111111101010010011001111;
         rom[22] = 24'b111111101011101111001100;
         rom[23] = 24'b111111010011010111011111;
         rom[24] = 24'b111111100100110101111010;
         rom[25] = 24'b111111011100100100000111;
         rom[26] = 24'b111111010000011000011110;
         rom[27] = 24'b111111010101101011110110;
         rom[28] = 24'b111111010010011111010001;
         rom[29] = 24'b111111100000110110011101;
         rom[30] = 24'b111111100011011110011001;
         rom[31] = 24'b111111101000011100110010;
         rom[32] = 24'b111111100111100000010010;
         rom[33] = 24'b111111101101111100010010;
         rom[34] = 24'b111111111010011110011110;
         rom[35] = 24'b111111101111111111100110;
         rom[36] = 24'b000000000101111111011000;
         rom[37] = 24'b000000000001001000010001;
         rom[38] = 24'b000000001110101111100000;
         rom[39] = 24'b000000001001100100001111;
         rom[40] = 24'b000000001011100101011110;
         rom[41] = 24'b000000011101100100010001;
         rom[42] = 24'b000000011011001011011010;
         rom[43] = 24'b000000011110001010100011;
         rom[44] = 24'b000000100100100001000010;
         rom[45] = 24'b000000101011011111100111;
         rom[46] = 24'b000000010110011111110011;
         rom[47] = 24'b000000100001011111000100;
         rom[48] = 24'b000000010000110110011110;
         rom[49] = 24'b000000101111000001111010;
         rom[50] = 24'b000000010100110001000010;
         rom[51] = 24'b000000010100110110010010;
         rom[52] = 24'b000000011010010010001111;
         rom[53] = 24'b000000000010000100111110;
         rom[54] = 24'b000000001110001001101101;
         rom[55] = 24'b111111111110000110111001;
         rom[56] = 24'b111111110111011111000010;
         rom[57] = 24'b111111110100110010100010;
         rom[58] = 24'b111111100101110000101011;
         rom[59] = 24'b111111110010110010101011;
         rom[60] = 24'b111111011100101100010100;
         rom[61] = 24'b111111011011011101000111;
         rom[62] = 24'b111111101000101010000011;
         rom[63] = 24'b111111010000001110111011;
         rom[64] = 24'b111111011000111001010010;
         rom[65] = 24'b111111100010100100111110;
         rom[66] = 24'b111111001110010111001010;
         rom[67] = 24'b111111011011100000100111;
         rom[68] = 24'b111111100101001011100011;
         rom[69] = 24'b111111101000111010100011;
         rom[70] = 24'b111111101000101001101001;
         rom[71] = 24'b000000000011000100111101;
         rom[72] = 24'b111111111001100011010111;
         rom[73] = 24'b000000000010110100101000;
         rom[74] = 24'b000000001011000101010000;
         rom[75] = 24'b000000010100011011000000;
         rom[76] = 24'b000000011010100100110100;
         rom[77] = 24'b000000011010100001000011;
         rom[78] = 24'b000000100101010011101011;
         rom[79] = 24'b000000100011111011010111;
         rom[80] = 24'b000000011111001110011001;
         rom[81] = 24'b000000100001101011000110;
         rom[82] = 24'b000000011110100100011100;
         rom[83] = 24'b000000110011000110100010;
         rom[84] = 24'b000000100001110111111100;
         rom[85] = 24'b000000011101100010011011;
         rom[86] = 24'b000000011000010101111000;
         rom[87] = 24'b000000011001011010111011;
         rom[88] = 24'b000000010100010110000100;
         rom[89] = 24'b000000011011011100100010;
         rom[90] = 24'b000000000001110100001111;
         rom[91] = 24'b111111111100100101000011;
         rom[92] = 24'b111111111110111010001001;
         rom[93] = 24'b111111101100101100011011;
         rom[94] = 24'b111111110000001000010001;
         rom[95] = 24'b111111100100011111010000;
         rom[96] = 24'b111111101000100100011110;
         rom[97] = 24'b111111110101000110001100;
         rom[98] = 24'b111111011010000111000001;
         rom[99] = 24'b111111011101101100010100;
         rom[100] = 24'b111111100001011010110110;
         rom[101] = 24'b111111011110010010111111;
         rom[102] = 24'b111111010010001010100110;
         rom[103] = 24'b111111010101001100000011;
         rom[104] = 24'b111111100101100000101001;
         rom[105] = 24'b111111100001100000111110;
         rom[106] = 24'b111111101011101101111110;
         rom[107] = 24'b111111110010001011000000;
         rom[108] = 24'b000000001001011001011111;
         rom[109] = 24'b000000010100001001111101;
         rom[110] = 24'b000000000000010110111101;
         rom[111] = 24'b111111111011000100011111;
         rom[112] = 24'b000000011011100100101001;
         rom[113] = 24'b000000000101011001011010;
         rom[114] = 24'b000000010011110010101011;
         rom[115] = 24'b000000100001001001010001;
         rom[116] = 24'b000000010101000110000001;
         rom[117] = 24'b000000101101111000011000;
         rom[118] = 24'b000000011010111001011101;
         rom[119] = 24'b000000100100111101111010;
         rom[120] = 24'b000000100101100110111111;
         rom[121] = 24'b000000001100011011000001;
         rom[122] = 24'b000000010010111010100001;
         rom[123] = 24'b000000001101110110001000;
         rom[124] = 24'b000000010001101001001101;
         rom[125] = 24'b000000001011100111100010;
         rom[126] = 24'b111111111111010111111011;
         rom[127] = 24'b111111111111101100101011;
         rom[128] = 24'b111111101100111111100010;
         rom[129] = 24'b111111110001010000001101;
         rom[130] = 24'b111111110010111010110101;
         rom[131] = 24'b111111110000111101011111;
         rom[132] = 24'b111111100010000100110001;
         rom[133] = 24'b111111101011011101010111;
         rom[134] = 24'b111111011010001101110000;
         rom[135] = 24'b111111100001011111110101;
         rom[136] = 24'b111111011011101111010001;
         rom[137] = 24'b111111011001001000001111;
         rom[138] = 24'b111111100001101100111110;
         rom[139] = 24'b111111011111111100001101;
         rom[140] = 24'b111111101001001011100001;
         rom[141] = 24'b111111110011100010011010;
         rom[142] = 24'b111111011100011011111011;
         rom[143] = 24'b111111111101011110011111;
         rom[144] = 24'b111111110110100101101110;
         rom[145] = 24'b111111111110000011010100;
         rom[146] = 24'b111111111101010011000111;
         rom[147] = 24'b000000000101101001010000;
         rom[148] = 24'b000000010100001110100110;
         rom[149] = 24'b000000010000011100100111;
         rom[150] = 24'b000000010111101111001011;
         rom[151] = 24'b000000011110101111001100;
         rom[152] = 24'b000000001111001011000110;
         rom[153] = 24'b000000101011100001001000;
         rom[154] = 24'b000000101001000000111000;
         rom[155] = 24'b000000011011111001100110;
         rom[156] = 24'b000000001110100111001001;
         rom[157] = 24'b000000100110011000011110;
         rom[158] = 24'b000000010110001101110100;
         rom[159] = 24'b000000010111100010111001;
         rom[160] = 24'b000000010010010010111000;
         rom[161] = 24'b000000000000110000000010;
         rom[162] = 24'b000000001000111010000011;
         rom[163] = 24'b000000000001101001010001;
         rom[164] = 24'b000000000010010111111110;
         rom[165] = 24'b111111110100011001001001;
         rom[166] = 24'b111111101110000011110110;
         rom[167] = 24'b111111101001000101111000;
         rom[168] = 24'b111111100000100101110011;
         rom[169] = 24'b111111100100011100100001;
         rom[170] = 24'b111111011110010010011101;
         rom[171] = 24'b111111010111011100100100;
         rom[172] = 24'b111111101100000010001000;
         rom[173] = 24'b111111011100111011011111;
         rom[174] = 24'b111111011000111001000001;
         rom[175] = 24'b111111100000000101100010;
         rom[176] = 24'b111111101011111110111011;
         rom[177] = 24'b111111011011001110010000;
         rom[178] = 24'b111111011010011100110011;
         rom[179] = 24'b111111110100000100111000;
         rom[180] = 24'b111111101111011010010000;
         rom[181] = 24'b000000000010011011100010;
         rom[182] = 24'b111111110100010011111101;
         rom[183] = 24'b000000000010010101110001;
         rom[184] = 24'b000000010010110100001101;
         rom[185] = 24'b000000001101100011001011;
         rom[186] = 24'b000000010011010001101010;
         rom[187] = 24'b000000011001001000110100;
         rom[188] = 24'b000000100111011100001111;
         rom[189] = 24'b000000011110001010000101;
         rom[190] = 24'b000000011110001011011111;
         rom[191] = 24'b000000100001110100000001;
         rom[192] = 24'b000000100011111111011111;
         rom[193] = 24'b000000100000010000011010;
         rom[194] = 24'b000000100101010000111100;
         rom[195] = 24'b000000011000111010010110;
         rom[196] = 24'b000000010111100000110100;
         rom[197] = 24'b000000001110101010100111;
         rom[198] = 24'b000000010011110010110010;
         rom[199] = 24'b000000001101101111110001;
         rom[200] = 24'b000000001001100101101011;
         rom[201] = 24'b111111110101100011101000;
         rom[202] = 24'b111111110000100110001010;
         rom[203] = 24'b111111111101100100010011;
         rom[204] = 24'b111111100010100011011111;
         rom[205] = 24'b111111011001000111111100;
         rom[206] = 24'b111111011100110100001101;
         rom[207] = 24'b111111100011110011100110;
         rom[208] = 24'b111111010000001110010100;
         rom[209] = 24'b111111011100001100010010;
         rom[210] = 24'b111111010111000111110011;
         rom[211] = 24'b111111100110011000010100;
         rom[212] = 24'b111111011010100011101000;
         rom[213] = 24'b111111010111010110101111;
         rom[214] = 24'b111111101110100110110110;
         rom[215] = 24'b111111111011101101100000;
         rom[216] = 24'b111111101110101100110100;
         rom[217] = 24'b111111110010000101111001;
         rom[218] = 24'b000000001001100010100110;
         rom[219] = 24'b111111111001110111010010;
         rom[220] = 24'b000000010100001000000010;
         rom[221] = 24'b000000001000010011111101;
         rom[222] = 24'b000000101001101101001001;
         rom[223] = 24'b000000001111000101111000;
         rom[224] = 24'b000000100000010100100000;
         rom[225] = 24'b000000100000000011000101;
         rom[226] = 24'b000000100000000000101001;
         rom[227] = 24'b000000100010100001001101;
         rom[228] = 24'b000000101011100100111110;
         rom[229] = 24'b000000011110111101111100;
         rom[230] = 24'b000000100110011010110110;
         rom[231] = 24'b000000100111100001000000;
         rom[232] = 24'b000000011001110001001010;
         rom[233] = 24'b000000010101100101100001;
         rom[234] = 24'b000000001001001111001000;
         rom[235] = 24'b000000001011001001011100;
         rom[236] = 24'b111111111010000011011000;
         rom[237] = 24'b000000000100001011110001;
         rom[238] = 24'b111111101101111011110011;
         rom[239] = 24'b111111101001101000110111;
         rom[240] = 24'b111111110000000001101100;
         rom[241] = 24'b111111100101010001100010;
         rom[242] = 24'b111111100000001101101011;
         rom[243] = 24'b111111100000110100110101;
         rom[244] = 24'b111111011101011010000110;
         rom[245] = 24'b111111010010010000111110;
         rom[246] = 24'b111111100111110000011100;
         rom[247] = 24'b111111010001010000011001;
         rom[248] = 24'b111111100011101010101011;
         rom[249] = 24'b111111100110111000000111;
         rom[250] = 24'b111111100101010001011110;
         rom[251] = 24'b111111101000011101110100;
         rom[252] = 24'b111111101011011111110111;
         rom[253] = 24'b111111100000110100001011;
         rom[254] = 24'b000000001000011010110111;
         rom[255] = 24'b000000000110100100010001;
         rom[256] = 24'b000000001111101000110011;
         rom[257] = 24'b000000001000001101110001;
         rom[258] = 24'b000000100011111110011000;
         rom[259] = 24'b000000100011010111000111;
         rom[260] = 24'b000000100111010100101001;
         rom[261] = 24'b000000100000101001100101;
         rom[262] = 24'b000000100001111101101001;
         rom[263] = 24'b000000101010011010000010;
         rom[264] = 24'b000000100001100000010101;
         rom[265] = 24'b000000100011000000100110;
         rom[266] = 24'b000000011011101111001111;
         rom[267] = 24'b000000010111101100000110;
         rom[268] = 24'b000000010100111001100100;
         rom[269] = 24'b000000010111111011110100;
         rom[270] = 24'b000000011000000010001001;
         rom[271] = 24'b000000001111001010111101;
         rom[272] = 24'b000000001000011101110100;
         rom[273] = 24'b111111110100110000000001;
         rom[274] = 24'b111111111101000010110001;
         rom[275] = 24'b111111110011111011011001;
         rom[276] = 24'b111111110111110111101011;
         rom[277] = 24'b111111100011111000101110;
         rom[278] = 24'b111111110100101011100001;
         rom[279] = 24'b111111101110010101011111;
         rom[280] = 24'b111111011111011101010100;
         rom[281] = 24'b111111011000101110101100;
         rom[282] = 24'b111111100011101100111000;
         rom[283] = 24'b111111011111000000101100;
         rom[284] = 24'b111111010011110011101000;
         rom[285] = 24'b111111100000111100110111;
         rom[286] = 24'b111111101110110000110001;
         rom[287] = 24'b111111100100001101100011;
         rom[288] = 24'b111111111000101010011000;
         rom[289] = 24'b111111111000011000010010;
         rom[290] = 24'b000000001001110111110011;
         rom[291] = 24'b111111111100100011100101;
         rom[292] = 24'b000000001101110011010101;
         rom[293] = 24'b000000001101110111111100;
         rom[294] = 24'b000000000001011111101011;
         rom[295] = 24'b000000011001000110000101;
         rom[296] = 24'b000000011111101011010011;
         rom[297] = 24'b000000100011111100100011;
         rom[298] = 24'b000000100101000000011110;
         rom[299] = 24'b000000100011111111001010;
         rom[300] = 24'b000000100100101011010111;
         rom[301] = 24'b000000100110000001000101;
         rom[302] = 24'b000000100000010001110001;
         rom[303] = 24'b000000100100111101001111;
         rom[304] = 24'b000000011001010110110100;
         rom[305] = 24'b000000011000011100010100;
         rom[306] = 24'b000000011000010110011101;
         rom[307] = 24'b000000000110010111000011;
         rom[308] = 24'b000000000111110000001100;
         rom[309] = 24'b111111101101011001011000;
         rom[310] = 24'b111111110111000001010001;
         rom[311] = 24'b111111101111011010100110;
         rom[312] = 24'b111111101110000000001000;
         rom[313] = 24'b111111100100001001101111;
         rom[314] = 24'b111111100010000110000011;
         rom[315] = 24'b111111011101000000100011;
         rom[316] = 24'b111111011101000101100000;
         rom[317] = 24'b111111101011010111111001;
         rom[318] = 24'b111111011000010101001001;
         rom[319] = 24'b111111100011000110010101;
         rom[320] = 24'b111111010101000000001110;
         rom[321] = 24'b111111101000110000100100;
         rom[322] = 24'b111111011001111101000010;
         rom[323] = 24'b111111101101110101001111;
         rom[324] = 24'b111111100110000011000100;
         rom[325] = 24'b111111101111100001111000;
         rom[326] = 24'b111111110111011001111110;
         rom[327] = 24'b111111111110110011110101;
         rom[328] = 24'b111111111000111111101011;
         rom[329] = 24'b000000001110101000010010;
         rom[330] = 24'b000000011000101001110101;
         rom[331] = 24'b000000010001000001101110;
         rom[332] = 24'b000000010101110100010111;
         rom[333] = 24'b000000100011110010101101;
         rom[334] = 24'b000000100100100010101001;
         rom[335] = 24'b000000100001011101001011;
         rom[336] = 24'b000000100011010010110101;
         rom[337] = 24'b000000110010001001001001;
         rom[338] = 24'b000000011101001001011000;
         rom[339] = 24'b000000100001111111111111;
         rom[340] = 24'b000000011110101000011101;
         rom[341] = 24'b000000011101111101000010;
         rom[342] = 24'b000000011111100100011110;
         rom[343] = 24'b000000001010100000100100;
         rom[344] = 24'b000000000100010110110101;
         rom[345] = 24'b111111111001010101000111;
         rom[346] = 24'b111111110010000110001111;
         rom[347] = 24'b111111101101100011111101;
         rom[348] = 24'b111111101100000001000010;
         rom[349] = 24'b111111101001101010010000;
         rom[350] = 24'b111111101101011010010011;
         rom[351] = 24'b111111010110110011000000;
         rom[352] = 24'b111111100100010010111111;
         rom[353] = 24'b111111100011001100111011;
         rom[354] = 24'b111111011010110101011111;
         rom[355] = 24'b111111010111001010111100;
         rom[356] = 24'b111111100100001100000111;
         rom[357] = 24'b111111011000110111100101;
         rom[358] = 24'b111111100110100111010110;
         rom[359] = 24'b111111100011110001001100;
         rom[360] = 24'b111111101000010010000110;
         rom[361] = 24'b111111101100010000110000;
         rom[362] = 24'b111111101011101001101011;
         rom[363] = 24'b111111111101001111000001;
         rom[364] = 24'b000000001001011010111001;
         rom[365] = 24'b000000001110100111110100;
         rom[366] = 24'b000000001101110010001010;
         rom[367] = 24'b000000011100101101111100;
         rom[368] = 24'b000000000111001110100001;
         rom[369] = 24'b000000011010011100010101;
         rom[370] = 24'b000000011101101100000010;
         rom[371] = 24'b000000110011000011000111;
         rom[372] = 24'b000000100101111110110000;
         rom[373] = 24'b000000011010101011110001;
         rom[374] = 24'b000000100111101000101111;
         rom[375] = 24'b000000100101110110101100;
         rom[376] = 24'b000000011000110010011011;
         rom[377] = 24'b000000100011100011111100;
         rom[378] = 24'b000000010111100011010101;
         rom[379] = 24'b000000010111000010100110;
         rom[380] = 24'b000000001011010000111011;
         rom[381] = 24'b000000010000100111101011;
         rom[382] = 24'b000000000010011000111111;
         rom[383] = 24'b111111110111110001000111;
         rom[384] = 24'b111111101111110011110111;
         rom[385] = 24'b111111101111101000011101;
         rom[386] = 24'b111111101011011100110011;
         rom[387] = 24'b111111011001010010011011;
         rom[388] = 24'b111111100100011011010101;
         rom[389] = 24'b111111011101101101100110;
         rom[390] = 24'b111111100001111101000111;
         rom[391] = 24'b111111011011100001011101;
         rom[392] = 24'b111111100010111000000110;
         rom[393] = 24'b111111100011010100010001;
         rom[394] = 24'b111111101001010001100100;
         rom[395] = 24'b111111100001100010011111;
         rom[396] = 24'b111111110111011111101111;
         rom[397] = 24'b111111100101110001000110;
         rom[398] = 24'b111111111110011101101110;
         rom[399] = 24'b000000000010111100100000;
         rom[400] = 24'b000000000001000101110011;
         rom[401] = 24'b000000000001000111101001;
         rom[402] = 24'b000000010010111100010001;
         rom[403] = 24'b000000000001001011011100;
         rom[404] = 24'b000000100001100000010011;
         rom[405] = 24'b000000011111111100111011;
         rom[406] = 24'b000000010101010000111110;
         rom[407] = 24'b000000100110000011110111;
         rom[408] = 24'b000000101101001001011100;
         rom[409] = 24'b000000010011001111110100;
         rom[410] = 24'b000000100111000011111011;
         rom[411] = 24'b000000011110011101011111;
         rom[412] = 24'b000000100010011001000101;
         rom[413] = 24'b000000100000001111100010;
         rom[414] = 24'b000000010011011111000011;
         rom[415] = 24'b000000010000100100001011;
         rom[416] = 24'b000000001010100110110100;
         rom[417] = 24'b111111111111001011011100;
         rom[418] = 24'b000000001010010100011101;
         rom[419] = 24'b111111100111111100100101;
         rom[420] = 24'b111111101100101100100001;
         rom[421] = 24'b111111101011100100111001;
         rom[422] = 24'b111111110010100011000010;
         rom[423] = 24'b111111100011111001001111;
         rom[424] = 24'b111111100001100111011101;
         rom[425] = 24'b111111011111010110001000;
         rom[426] = 24'b111111010110000001111110;
         rom[427] = 24'b111111011101010100000100;
         rom[428] = 24'b111111100010000011010010;
         rom[429] = 24'b111111011110110110001100;
         rom[430] = 24'b111111010000001001110011;
         rom[431] = 24'b111111100000111101110111;
         rom[432] = 24'b111111100011100000001100;
         rom[433] = 24'b111111110001011101101111;
         rom[434] = 24'b111111101100001011010100;
         rom[435] = 24'b111111111001001110000101;
         rom[436] = 24'b111111111001110100111100;
         rom[437] = 24'b111111111001000011000001;
         rom[438] = 24'b000000001011010100011001;
         rom[439] = 24'b000000010110111001110011;
         rom[440] = 24'b000000011001011100110000;
         rom[441] = 24'b000000011000000100000111;
         rom[442] = 24'b000000011001110011100100;
         rom[443] = 24'b000000010000011110001111;
         rom[444] = 24'b000000100110111111010010;
         rom[445] = 24'b000000100000100011001111;
         rom[446] = 24'b000000011001011111111110;
         rom[447] = 24'b000000100011101100001110;
         rom[448] = 24'b000000100010000101001011;
         rom[449] = 24'b000000101011101111001100;
         rom[450] = 24'b000000001110011001001011;
         rom[451] = 24'b000000011001111000111001;
         rom[452] = 24'b000000010001011001000011;
         rom[453] = 24'b000000001110001111010000;
         rom[454] = 24'b000000001001001100111111;
         rom[455] = 24'b000000001000011000101100;
         rom[456] = 24'b111111101000011011000111;
         rom[457] = 24'b111111100111001110110010;
         rom[458] = 24'b111111100111001101111011;
         rom[459] = 24'b111111011011011111110101;
         rom[460] = 24'b111111010011111100110000;
         rom[461] = 24'b111111100001110011011111;
         rom[462] = 24'b111111100111011110101010;
         rom[463] = 24'b111111011110000000101111;
         rom[464] = 24'b111111001011000101001111;
         rom[465] = 24'b111111010101100000011010;
         rom[466] = 24'b111111011110001001100000;
         rom[467] = 24'b111111010101010010100001;
         rom[468] = 24'b111111110000100011100010;
         rom[469] = 24'b111111101101000000111110;
         rom[470] = 24'b111111110000111111100111;
         rom[471] = 24'b111111110011010110100101;
         rom[472] = 24'b000000000001010011001101;
         rom[473] = 24'b000000000100100111111100;
         rom[474] = 24'b000000000011010100111101;
         rom[475] = 24'b000000001011111101010001;
         rom[476] = 24'b000000100011110010110111;
         rom[477] = 24'b000000010001010001110100;
         rom[478] = 24'b000000100001111110101111;
         rom[479] = 24'b000000101110100001101100;
         rom[480] = 24'b000000011111110011000000;
         rom[481] = 24'b000000101001110010010110;
         rom[482] = 24'b000000110111111010111111;
         rom[483] = 24'b000000011010111001110101;
         rom[484] = 24'b000000011100011110001010;
         rom[485] = 24'b000000101011000010010011;
         rom[486] = 24'b000000100110011001101101;
         rom[487] = 24'b000000010101001100001110;
         rom[488] = 24'b000000001111100001000000;
         rom[489] = 24'b111111111111110001011010;
         rom[490] = 24'b000000001011111100110011;
         rom[491] = 24'b000000001100011101110001;
         rom[492] = 24'b111111111011001000000001;
         rom[493] = 24'b111111101100110000100001;
         rom[494] = 24'b111111101100001110101100;
         rom[495] = 24'b111111100010100110101100;
         rom[496] = 24'b111111100011101000001101;
         rom[497] = 24'b111111100000101100000111;
         rom[498] = 24'b111111100001111101101100;
         rom[499] = 24'b111111001110110100000011;
         rom[500] = 24'b111111100101011111010011;
         rom[501] = 24'b111111011010111101110111;
         rom[502] = 24'b111111011000100001101100;
         rom[503] = 24'b111111100001110011010011;
         rom[504] = 24'b111111011101111101001110;
         rom[505] = 24'b111111100011111000011110;
         rom[506] = 24'b111111101001111100001100;
         rom[507] = 24'b111111100111101001101111;
         rom[508] = 24'b111111110101011111111000;
         rom[509] = 24'b000000000110111111111000;
         rom[510] = 24'b000000010001101011101010;
         rom[511] = 24'b000000001011110110101010;
         rom[512] = 24'b000000010110101010110000;
         rom[513] = 24'b000000010110101100110110;
         rom[514] = 24'b000000001111000110110010;
         rom[515] = 24'b000000011110011110100000;
         rom[516] = 24'b000000101100101011000111;
         rom[517] = 24'b000000100110000000011100;
         rom[518] = 24'b000000101000000001001010;
         rom[519] = 24'b000000011101110101011000;
         rom[520] = 24'b000000010110110001100010;
         rom[521] = 24'b000000100000001010000010;
         rom[522] = 24'b000000011011001100011011;
         rom[523] = 24'b000000001101001001011010;
         rom[524] = 24'b000000000111001010110101;
         rom[525] = 24'b000000001001100000101110;
         rom[526] = 24'b000000001010110001001000;
         rom[527] = 24'b000000000100001010010011;
         rom[528] = 24'b000000000011010000001001;
         rom[529] = 24'b111111101101011010001011;
         rom[530] = 24'b111111101110011000011100;
         rom[531] = 24'b111111011110110101011100;
         rom[532] = 24'b111111100011001111000000;
         rom[533] = 24'b111111010100010100001010;
         rom[534] = 24'b111111101001010010001011;
         rom[535] = 24'b111111011001010101111100;
         rom[536] = 24'b111111011001010011000111;
         rom[537] = 24'b111111100001100100111001;
         rom[538] = 24'b111111010111111110000011;
         rom[539] = 24'b111111011101100110101111;
         rom[540] = 24'b111111100000001100000111;
         rom[541] = 24'b111111100111011101110011;
         rom[542] = 24'b111111101010000000110110;
         rom[543] = 24'b000000000000110110010010;
         rom[544] = 24'b111111110101011101001101;
         rom[545] = 24'b111111111110111001100110;
         rom[546] = 24'b000000001000001100011100;
         rom[547] = 24'b000000000111111001010001;
         rom[548] = 24'b000000011010000111101110;
         rom[549] = 24'b000000010001000110101001;
         rom[550] = 24'b000000001000101010101110;
         rom[551] = 24'b000000011110110110001011;
         rom[552] = 24'b000000011110010111110001;
         rom[553] = 24'b000000100010100100010000;
         rom[554] = 24'b000000110010110000010000;
         rom[555] = 24'b000000101010011110110010;
         rom[556] = 24'b000000100100000101101110;
         rom[557] = 24'b000000101100010110000000;
         rom[558] = 24'b000000011011010001000010;
         rom[559] = 24'b000000011100001100010100;
         rom[560] = 24'b000000010100110110000111;
         rom[561] = 24'b000000100001010101000001;
         rom[562] = 24'b000000001110101110001101;
         rom[563] = 24'b000000000101001101100010;
         rom[564] = 24'b111111110011000111110011;
         rom[565] = 24'b111111110101010100110001;
         rom[566] = 24'b111111101000010110010100;
         rom[567] = 24'b111111110011000010001001;
         rom[568] = 24'b111111100100000010011110;
         rom[569] = 24'b111111010101001110000100;
         rom[570] = 24'b111111010111101011110111;
         rom[571] = 24'b111111100000011101111000;
         rom[572] = 24'b111111010110101101101111;
         rom[573] = 24'b111111011101111010010110;
         rom[574] = 24'b111111101010010000011010;
         rom[575] = 24'b111111100100111110101111;
         rom[576] = 24'b111111101111010110100001;
         rom[577] = 24'b111111100000101111101100;
         rom[578] = 24'b111111101100011110000100;
         rom[579] = 24'b111111101000000101100100;
         rom[580] = 24'b111111110011101000011010;
         rom[581] = 24'b111111111011111100100001;
         rom[582] = 24'b111111111110111000100011;
         rom[583] = 24'b000000010001000001010000;
         rom[584] = 24'b000000011001010000101111;
         rom[585] = 24'b000000010101100111011111;
         rom[586] = 24'b000000010101010001110001;
         rom[587] = 24'b000000011011100101000010;
         rom[588] = 24'b000000011001000110111111;
         rom[589] = 24'b000000100000010100110111;
         rom[590] = 24'b000000100001100111101101;
         rom[591] = 24'b000000101110010110010111;
         rom[592] = 24'b000000100000100000000110;
         rom[593] = 24'b000000011111110000110010;
         rom[594] = 24'b000000101010111010100111;
         rom[595] = 24'b000000010001000101001110;
         rom[596] = 24'b000000010100101011010010;
         rom[597] = 24'b000000010100001100011100;
         rom[598] = 24'b000000000111110110011011;
         rom[599] = 24'b000000001111001011000001;
         rom[600] = 24'b111111111001110110110110;
         rom[601] = 24'b111111110111010010010001;
         rom[602] = 24'b111111100101101010000001;
         rom[603] = 24'b111111101100100111101111;
         rom[604] = 24'b111111110011000111111011;
         rom[605] = 24'b111111100010001011011011;
         rom[606] = 24'b111111101110010110111101;
         rom[607] = 24'b111111011100100110011001;
         rom[608] = 24'b111111001110001001111001;
         rom[609] = 24'b111111011100011010010010;
         rom[610] = 24'b111111100000111101011010;
         rom[611] = 24'b111111011101101010011111;
         rom[612] = 24'b111111011111100110101011;
         rom[613] = 24'b111111100010010010110110;
         rom[614] = 24'b111111110011100100101100;
         rom[615] = 24'b111111101101101011010011;
         rom[616] = 24'b111111110010000111011000;
         rom[617] = 24'b000000000110100001100100;
         rom[618] = 24'b111111110111100001001000;
         rom[619] = 24'b111111111001010000001110;
         rom[620] = 24'b000000010001001101000001;
         rom[621] = 24'b000000010001011010011011;
         rom[622] = 24'b000000011000110000001100;
         rom[623] = 24'b000000011100011001100111;
         rom[624] = 24'b000000011110001100010110;
         rom[625] = 24'b000000100001001111010100;
         rom[626] = 24'b000000010011110001111001;
         rom[627] = 24'b000000011001011010101110;
         rom[628] = 24'b000000101000000100011000;
         rom[629] = 24'b000000101101101101010010;
         rom[630] = 24'b000000010111011010100001;
         rom[631] = 24'b000000010010001010110101;
         rom[632] = 24'b000000100000111111000001;
         rom[633] = 24'b000000010100000110010110;
         rom[634] = 24'b000000001011110001010001;
         rom[635] = 24'b000000001001001010011000;
         rom[636] = 24'b000000001001001100011011;
         rom[637] = 24'b111111111010011110101010;
         rom[638] = 24'b111111101101011111110000;
         rom[639] = 24'b111111111100001100001111;
         rom[640] = 24'b111111100110000010100100;
         rom[641] = 24'b111111011100010110101011;
         rom[642] = 24'b111111011110110000110111;
         rom[643] = 24'b111111100011110110111111;
         rom[644] = 24'b111111010101001100100100;
         rom[645] = 24'b111111011011011101100010;
         rom[646] = 24'b111111011011111101010000;
         rom[647] = 24'b111111011111010000110000;
         rom[648] = 24'b111111011000010001111110;
         rom[649] = 24'b111111011110100001001010;
         rom[650] = 24'b111111011111111101001110;
         rom[651] = 24'b111111101011011100001010;
         rom[652] = 24'b111111111101001100111111;
         rom[653] = 24'b111111111101111111000010;
         rom[654] = 24'b000000001110010000101010;
         rom[655] = 24'b000000000011010101000011;
         rom[656] = 24'b000000001001111110111000;
         rom[657] = 24'b000000001100000100111011;
         rom[658] = 24'b000000010001110111011111;
         rom[659] = 24'b000000011001110101110000;
         rom[660] = 24'b000000011110100000010000;
         rom[661] = 24'b000000011100000110001000;
         rom[662] = 24'b000000100101000111101100;
         rom[663] = 24'b000000100111011010010111;
         rom[664] = 24'b000000100111001001011101;
         rom[665] = 24'b000000100011000010100000;
         rom[666] = 24'b000000101001011001101111;
         rom[667] = 24'b000000011110010111001001;
         rom[668] = 24'b000000011010000000101110;
         rom[669] = 24'b000000001010000100010111;
         rom[670] = 24'b000000001110010010010110;
         rom[671] = 24'b000000011010001100011101;
         rom[672] = 24'b000000001100101110011001;
         rom[673] = 24'b111111101101110111111100;
         rom[674] = 24'b000000000001010100001010;
         rom[675] = 24'b111111110110111111111000;
         rom[676] = 24'b111111100100010111111000;
         rom[677] = 24'b111111101000110000111001;
         rom[678] = 24'b111111100101000110010110;
         rom[679] = 24'b111111101011110001111001;
         rom[680] = 24'b111111011000110000101010;
         rom[681] = 24'b111111010011110001000101;
         rom[682] = 24'b111111011111111001011001;
         rom[683] = 24'b111111100010100010101111;
         rom[684] = 24'b111111011010010011100101;
         rom[685] = 24'b111111101010011000100110;
         rom[686] = 24'b111111100001111011101101;
         rom[687] = 24'b111111100111101000110111;
         rom[688] = 24'b111111100100101001010011;
         rom[689] = 24'b111111111011110001010001;
         rom[690] = 24'b000000000001000111110110;
         rom[691] = 24'b000000000001110011111100;
         rom[692] = 24'b111111111000101101110110;
         rom[693] = 24'b000000010101010010111100;
         rom[694] = 24'b000000011000001001100001;
         rom[695] = 24'b000000010110000011101001;
         rom[696] = 24'b000000010111001110011111;
         rom[697] = 24'b000000011001101110001001;
         rom[698] = 24'b000000010111001111110011;
         rom[699] = 24'b000000010110100001110101;
         rom[700] = 24'b000000100100001110011011;
         rom[701] = 24'b000000011101111001000001;
         rom[702] = 24'b000000100101010010010011;
         rom[703] = 24'b000000100011001010100010;
         rom[704] = 24'b000000011001100010110011;
         rom[705] = 24'b000000011001000110100010;
         rom[706] = 24'b000000011000011110010101;
         rom[707] = 24'b000000001110001011001110;
         rom[708] = 24'b000000001111110100000100;
         rom[709] = 24'b000000000000110101010111;
         rom[710] = 24'b111111110110000000111100;
         rom[711] = 24'b111111101011111101111110;
         rom[712] = 24'b111111100011001111101011;
         rom[713] = 24'b111111101110001110001100;
         rom[714] = 24'b111111101101110111101110;
         rom[715] = 24'b111111101100010011011111;
         rom[716] = 24'b111111011000111011111011;
         rom[717] = 24'b111111100001010111101000;
         rom[718] = 24'b111111010100001111111100;
         rom[719] = 24'b111111100010010101000111;
         rom[720] = 24'b111111011010100001010001;
         rom[721] = 24'b111111101110111011010010;
         rom[722] = 24'b111111101000011010101101;
         rom[723] = 24'b111111100011000000100101;
         rom[724] = 24'b111111111000111011111110;
         rom[725] = 24'b111111110110110001101111;
         rom[726] = 24'b000000000010000001011101;
         rom[727] = 24'b111111111010101000100001;
         rom[728] = 24'b000000001101001110001100;
         rom[729] = 24'b000000010111011100111100;
         rom[730] = 24'b000000001100101011110000;
         rom[731] = 24'b000000010000001101100101;
         rom[732] = 24'b000000100011011111110000;
         rom[733] = 24'b000000011010001101010000;
         rom[734] = 24'b000000100100010001010100;
         rom[735] = 24'b000000011111010010101111;
         rom[736] = 24'b000000100110010000010101;
         rom[737] = 24'b000000101000011001001111;
         rom[738] = 24'b000000100111110110100111;
         rom[739] = 24'b000000010010110011011011;
         rom[740] = 24'b000000010011010101110010;
         rom[741] = 24'b000000001111110001100010;
         rom[742] = 24'b000000011001101100101110;
         rom[743] = 24'b000000010100101101111010;
         rom[744] = 24'b000000000101011100101000;
         rom[745] = 24'b000000000111010110111100;
         rom[746] = 24'b000000000110110001100101;
         rom[747] = 24'b111111110100110101001111;
         rom[748] = 24'b111111101111111110101000;
         rom[749] = 24'b111111101001110111010101;
         rom[750] = 24'b111111011100011001101101;
         rom[751] = 24'b111111100101100110101001;
         rom[752] = 24'b111111001110110010110010;
         rom[753] = 24'b111111100111101000111011;
         rom[754] = 24'b111111100111010110011110;
         rom[755] = 24'b111111100000111101011110;
         rom[756] = 24'b111111100010001110011111;
         rom[757] = 24'b111111100000111010000000;
         rom[758] = 24'b111111110011110000000010;
         rom[759] = 24'b111111100011110000101100;
         rom[760] = 24'b111111100001100011111101;
         rom[761] = 24'b111111111011111000101101;
         rom[762] = 24'b111111110000110000001100;
         rom[763] = 24'b000000000010101010110101;
         rom[764] = 24'b111111110111100111011001;
         rom[765] = 24'b111111111111110011111001;
         rom[766] = 24'b000000010101111010110111;
         rom[767] = 24'b000000010010111111010001;
         rom[768] = 24'b000000011111100111011010;
         rom[769] = 24'b000000011110000110101101;
         rom[770] = 24'b000000101001010001010001;
         rom[771] = 24'b000000110001101010111111;
         rom[772] = 24'b000000011100010101101101;
         rom[773] = 24'b000000101010100110110011;
         rom[774] = 24'b000000011111101100100100;
         rom[775] = 24'b000000100100101010011101;
         rom[776] = 24'b000000011100101010110111;
         rom[777] = 24'b000000011110100010011011;
         rom[778] = 24'b000000011001010010101000;
         rom[779] = 24'b000000010011101100100110;
         rom[780] = 24'b000000000001011101011101;
         rom[781] = 24'b111111111001111000110101;
         rom[782] = 24'b000000000111001010001011;
         rom[783] = 24'b111111111010110001101100;
         rom[784] = 24'b111111101111011100110110;
         rom[785] = 24'b111111111011111000010101;
         rom[786] = 24'b111111101100100111011111;
         rom[787] = 24'b111111110000000011111001;
         rom[788] = 24'b111111100001110011001000;
         rom[789] = 24'b111111011100111101001110;
         rom[790] = 24'b111111011100001001111011;
         rom[791] = 24'b111111010010101100000000;
         rom[792] = 24'b111111100001011111110110;
         rom[793] = 24'b111111011110000101010011;
         rom[794] = 24'b111111100001001001011101;
         rom[795] = 24'b111111110011001010010110;
         rom[796] = 24'b111111110011111110100100;
         rom[797] = 24'b111111110001111100011010;
         rom[798] = 24'b111111110101000101100101;
         rom[799] = 24'b000000000110101010110001;
         rom[800] = 24'b111111111011011000101001;
         rom[801] = 24'b000000001000101111010000;
         rom[802] = 24'b000000000011111000101001;
         rom[803] = 24'b000000011100101110000111;
         rom[804] = 24'b000000100001001110001010;
         rom[805] = 24'b000000010111111010000110;
         rom[806] = 24'b000000011001001001000000;
         rom[807] = 24'b000000100110101110100011;
         rom[808] = 24'b000000101011011101011100;
         rom[809] = 24'b000000100000111011111001;
         rom[810] = 24'b000000010111011111101100;
         rom[811] = 24'b000000100011111010001000;
         rom[812] = 24'b000000011100100101001101;
         rom[813] = 24'b000000010111010101011011;
         rom[814] = 24'b000000010010010101011001;
         rom[815] = 24'b000000010111001000100011;
         rom[816] = 24'b000000010010111110000100;
         rom[817] = 24'b000000000011000000000000;
         rom[818] = 24'b111111110111000000110110;
         rom[819] = 24'b111111110101001111000001;
         rom[820] = 24'b111111111000011001110011;
         rom[821] = 24'b111111101010000010111001;
         rom[822] = 24'b111111110010100111110100;
         rom[823] = 24'b111111100100100011011001;
         rom[824] = 24'b111111100110001001001101;
         rom[825] = 24'b111111011110000010111010;
         rom[826] = 24'b111111100000000000000100;
         rom[827] = 24'b111111001111000111001111;
         rom[828] = 24'b111111100011110001000110;
         rom[829] = 24'b111111011101101000011001;
         rom[830] = 24'b111111100100100101110111;
         rom[831] = 24'b111111011010100010101101;
         rom[832] = 24'b111111101100110000010111;
         rom[833] = 24'b111111110010011000000001;
         rom[834] = 24'b111111101010011000010111;
         rom[835] = 24'b111111110101111000111000;
         rom[836] = 24'b111111111101011101110100;
         rom[837] = 24'b000000000001010000010100;
         rom[838] = 24'b000000010101000110100101;
         rom[839] = 24'b000000010001011100100100;
         rom[840] = 24'b000000011011000110001011;
         rom[841] = 24'b000000010111001100100101;
         rom[842] = 24'b000000101010110110101000;
         rom[843] = 24'b000000100100001010001001;
         rom[844] = 24'b000000100011111010100001;
         rom[845] = 24'b000000100101000101011001;
         rom[846] = 24'b000000100110100000001001;
         rom[847] = 24'b000000011001001101011100;
         rom[848] = 24'b000000100110010110110100;
         rom[849] = 24'b000000010110011000100101;
         rom[850] = 24'b000000011010011010011010;
         rom[851] = 24'b000000011010010110010100;
         rom[852] = 24'b000000001011000101100000;
         rom[853] = 24'b000000001000001111101101;
         rom[854] = 24'b111111111011100001010111;
         rom[855] = 24'b111111111110100100001010;
         rom[856] = 24'b111111111111000010001010;
         rom[857] = 24'b111111110110010111011111;
         rom[858] = 24'b111111100111001101110001;
         rom[859] = 24'b111111100110011111110000;
         rom[860] = 24'b111111011111111011111010;
         rom[861] = 24'b111111011001010011000100;
         rom[862] = 24'b111111011111100000111101;
         rom[863] = 24'b111111100100111001011001;
         rom[864] = 24'b111111011010101011110100;
         rom[865] = 24'b111111010101100110000010;
         rom[866] = 24'b111111100001010110101011;
         rom[867] = 24'b111111100100100100001001;
         rom[868] = 24'b111111101010100000110101;
         rom[869] = 24'b111111100011111100111100;
         rom[870] = 24'b111111101111111110011001;
         rom[871] = 24'b111111101101010100000111;
         rom[872] = 24'b000000000011100101001100;
         rom[873] = 24'b111111111001000110010111;
         rom[874] = 24'b000000000011010111101111;
         rom[875] = 24'b000000001001001000110100;
         rom[876] = 24'b000000010100001100000110;
         rom[877] = 24'b000000011110101110000010;
         rom[878] = 24'b000000010101111101101000;
         rom[879] = 24'b000000101010101001001100;
         rom[880] = 24'b000000011000000011001001;
         rom[881] = 24'b000000100101110100011111;
         rom[882] = 24'b000000100111011111011100;
         rom[883] = 24'b000000100101111110001000;
         rom[884] = 24'b000000100011001010110010;
         rom[885] = 24'b000000100000001001011000;
         rom[886] = 24'b000000011101011101011101;
         rom[887] = 24'b000000010110110111110011;
         rom[888] = 24'b000000001100011100110101;
         rom[889] = 24'b000000010010110000000111;
         rom[890] = 24'b000000000000001111110000;
         rom[891] = 24'b000000000101101110010111;
         rom[892] = 24'b111111111011100001101000;
         rom[893] = 24'b111111111010011010110100;
         rom[894] = 24'b111111100110111100110100;
         rom[895] = 24'b111111101101101101100111;
         rom[896] = 24'b111111010111010111011111;
         rom[897] = 24'b111111011101010101000101;
         rom[898] = 24'b111111100110000111101000;
         rom[899] = 24'b111111101001110101010100;
         rom[900] = 24'b111111011001101101011001;
         rom[901] = 24'b111111011010001000000001;
         rom[902] = 24'b111111100000110001011111;
         rom[903] = 24'b111111011000011110111000;
         rom[904] = 24'b111111010101110110111110;
         rom[905] = 24'b111111101101011111000001;
         rom[906] = 24'b111111101001001000010110;
         rom[907] = 24'b111111101000110111001001;
         rom[908] = 24'b111111111000110110000011;
         rom[909] = 24'b000000000001011110110111;
         rom[910] = 24'b111111111110000100000010;
         rom[911] = 24'b000000000010101000000111;
         rom[912] = 24'b000000010111101100100110;
         rom[913] = 24'b000000011110001101010010;
         rom[914] = 24'b000000010011111111000101;
         rom[915] = 24'b000000100111110000010010;
         rom[916] = 24'b000000100000110111010011;
         rom[917] = 24'b000000101101110011001110;
         rom[918] = 24'b000000101010011011000110;
         rom[919] = 24'b000000101010110001110000;
         rom[920] = 24'b000000100100111110001111;
         rom[921] = 24'b000000010101101000101101;
         rom[922] = 24'b000000100000111010000011;
         rom[923] = 24'b000000100001101010001010;
         rom[924] = 24'b000000010100111111101011;
         rom[925] = 24'b000000001011111110011111;
         rom[926] = 24'b000000011001100110011100;
         rom[927] = 24'b000000000001111110011101;
         rom[928] = 24'b111111111000100111101000;
         rom[929] = 24'b111111111000011000001000;
         rom[930] = 24'b111111101001111001110001;
         rom[931] = 24'b111111101101000000100100;
         rom[932] = 24'b111111011101101111010110;
         rom[933] = 24'b111111100010000010100111;
         rom[934] = 24'b111111101000010010001011;
         rom[935] = 24'b111111100100010110111001;
         rom[936] = 24'b111111010110110110100111;
         rom[937] = 24'b111111011000111000011011;
         rom[938] = 24'b111111011111001011010100;
         rom[939] = 24'b111111100000110101110000;
         rom[940] = 24'b111111011100000001111010;
         rom[941] = 24'b111111100100010101011110;
         rom[942] = 24'b111111101000111100010111;
         rom[943] = 24'b111111101101100101101111;
         rom[944] = 24'b111111110101100111000000;
         rom[945] = 24'b111111111100111010100001;
         rom[946] = 24'b111111111110000111110110;
         rom[947] = 24'b000000000001101101011100;
         rom[948] = 24'b000000001110101001111110;
         rom[949] = 24'b000000011111001001011001;
         rom[950] = 24'b000000010101101010000110;
         rom[951] = 24'b000000011010100111110111;
         rom[952] = 24'b000000011010001111111000;
         rom[953] = 24'b000000100000110110110101;
         rom[954] = 24'b000000101000000001010011;
         rom[955] = 24'b000000100011001011101001;
         rom[956] = 24'b000000100111011100011101;
         rom[957] = 24'b000000101100010010110111;
         rom[958] = 24'b000000100001010011010110;
         rom[959] = 24'b000000100001111010101010;
         rom[960] = 24'b000000100001000010010000;
         rom[961] = 24'b000000001110010010001000;
         rom[962] = 24'b000000000010100100000111;
         rom[963] = 24'b000000001111000100111000;
         rom[964] = 24'b000000000101111111011000;
         rom[965] = 24'b111111111110010011011100;
         rom[966] = 24'b111111111011111110010010;
         rom[967] = 24'b111111100001000110000010;
         rom[968] = 24'b111111011101001100101001;
         rom[969] = 24'b111111100111001001100110;
         rom[970] = 24'b111111010101110010100000;
         rom[971] = 24'b111111101001010110000101;
         rom[972] = 24'b111111100010111101000111;
         rom[973] = 24'b111111100101110100001100;
         rom[974] = 24'b111111010001001001100110;
         rom[975] = 24'b111111011011110110101000;
         rom[976] = 24'b111111101001011001110001;
         rom[977] = 24'b111111100011010111100110;
         rom[978] = 24'b111111101000110101000001;
         rom[979] = 24'b111111100101011011001110;
         rom[980] = 24'b111111101110101110010011;
         rom[981] = 24'b000000000000011011100011;
         rom[982] = 24'b000000000100110110100101;
         rom[983] = 24'b000000000100110110011100;
         rom[984] = 24'b000000010000000011001010;
         rom[985] = 24'b000000010110010001100010;
         rom[986] = 24'b000000010111100010110011;
         rom[987] = 24'b000000011010111101011001;
         rom[988] = 24'b000000010101001001000000;
         rom[989] = 24'b000000010011101001101001;
         rom[990] = 24'b000000100011100010100100;
         rom[991] = 24'b000000101010000111110000;
         rom[992] = 24'b000000011000100011010111;
         rom[993] = 24'b000000010101011110101101;
         rom[994] = 24'b000000011010100000100111;
         rom[995] = 24'b000000010101000011111111;
         rom[996] = 24'b000000100001111001001110;
         rom[997] = 24'b000000001011001111100101;
         rom[998] = 24'b000000011000001100100010;
         rom[999] = 24'b000000010101000100110000;
         rom[1000] = 24'b000000001011110100011110;
         rom[1001] = 24'b000000000110100000110111;
         rom[1002] = 24'b111111101000000100011001;
         rom[1003] = 24'b111111100001110000000110;
         rom[1004] = 24'b111111100001111010101000;
         rom[1005] = 24'b111111011011101010110101;
         rom[1006] = 24'b111111100000110110110101;
         rom[1007] = 24'b111111011100101110011111;
         rom[1008] = 24'b111111011011111010111100;
         rom[1009] = 24'b111111011110101110001101;
         rom[1010] = 24'b111111010000000100000100;
         rom[1011] = 24'b111111011000011011101010;
         rom[1012] = 24'b111111100100011101000011;
         rom[1013] = 24'b111111101011000001001100;
         rom[1014] = 24'b111111101111001010000010;
         rom[1015] = 24'b111111110010010110010110;
         rom[1016] = 24'b111111111110111110000100;
         rom[1017] = 24'b000000000100001010111101;
         rom[1018] = 24'b111111110111100011111011;
         rom[1019] = 24'b000000000100001100000001;
         rom[1020] = 24'b000000000110011111011010;
         rom[1021] = 24'b000000000100000011101110;
         rom[1022] = 24'b000000001111011001100100;
         rom[1023] = 24'b000000010101001011011010;
         rom[1024] = 24'b000000011000110000001110;
         rom[1025] = 24'b000000100110100001000111;
         rom[1026] = 24'b000000101011011101000110;
         rom[1027] = 24'b000000110011000100100000;
         rom[1028] = 24'b000000101110110110010100;
         rom[1029] = 24'b000000101001000000100100;
         rom[1030] = 24'b000000101010110001010110;
         rom[1031] = 24'b000000010100100111111110;
         rom[1032] = 24'b000000010100110011011010;
         rom[1033] = 24'b000000010101110010000101;
         rom[1034] = 24'b000000000110000101111111;
         rom[1035] = 24'b000000001111100001000100;
         rom[1036] = 24'b111111111101100001101000;
         rom[1037] = 24'b000000000010110101010010;
         rom[1038] = 24'b111111110011011111010111;
         rom[1039] = 24'b111111110111010001101001;
         rom[1040] = 24'b111111100111111010101101;
         rom[1041] = 24'b111111100111010001100111;
         rom[1042] = 24'b111111100100000010110011;
         rom[1043] = 24'b111111100101010010001100;
         rom[1044] = 24'b111111100100100010101101;
         rom[1045] = 24'b111111011001100010111110;
         rom[1046] = 24'b111111011101010111010111;
         rom[1047] = 24'b111111011111110001110110;
         rom[1048] = 24'b111111100000110101010110;
         rom[1049] = 24'b111111100011101101000101;
         rom[1050] = 24'b111111100101000000110011;
         rom[1051] = 24'b111111100110000111111001;
         rom[1052] = 24'b111111110010010110000010;
         rom[1053] = 24'b111111110011010000101101;
         rom[1054] = 24'b111111111111001110011011;
         rom[1055] = 24'b000000010001110101111010;
         rom[1056] = 24'b000000001101110100100100;
         rom[1057] = 24'b000000011001000011110100;
         rom[1058] = 24'b000000100001011001111000;
         rom[1059] = 24'b000000010101100001001101;
         rom[1060] = 24'b000000100001111011011010;
         rom[1061] = 24'b000000100001100100001110;
         rom[1062] = 24'b000000101101100111100110;
         rom[1063] = 24'b000000101110111101100000;
         rom[1064] = 24'b000000100100001010100010;
         rom[1065] = 24'b000000100011101010101000;
         rom[1066] = 24'b000000011000001100110111;
         rom[1067] = 24'b000000010110111100110010;
         rom[1068] = 24'b000000010101111111111000;
         rom[1069] = 24'b000000010001100011110110;
         rom[1070] = 24'b000000010100001011000011;
         rom[1071] = 24'b000000001000010110101011;
         rom[1072] = 24'b111111111111000101111010;
         rom[1073] = 24'b111111111100001111110011;
         rom[1074] = 24'b111111111001100011100010;
         rom[1075] = 24'b111111110010000111010111;
         rom[1076] = 24'b111111110000110000111000;
         rom[1077] = 24'b111111100111001100111011;
         rom[1078] = 24'b111111100011100011011110;
         rom[1079] = 24'b111111101001100100010101;
         rom[1080] = 24'b111111010101111000000011;
         rom[1081] = 24'b111111100011100001000011;
         rom[1082] = 24'b111111101111010011101100;
         rom[1083] = 24'b111111010111010101010110;
         rom[1084] = 24'b111111110010110101110100;
         rom[1085] = 24'b111111100111111100001000;
         rom[1086] = 24'b111111011000111100101110;
         rom[1087] = 24'b111111010101001000000110;
         rom[1088] = 24'b111111101011000110101101;
         rom[1089] = 24'b111111100111011100001001;
         rom[1090] = 24'b000000000010000010001101;
         rom[1091] = 24'b111111111001100000010011;
         rom[1092] = 24'b000000010010000000101001;
         rom[1093] = 24'b000000011000100100110011;
         rom[1094] = 24'b000000001100110110000100;
         rom[1095] = 24'b000000010110001010010100;
         rom[1096] = 24'b000000001010011000010101;
         rom[1097] = 24'b000000100100011011101010;
         rom[1098] = 24'b000000100100110010010001;
         rom[1099] = 24'b000000100000100100011011;
         rom[1100] = 24'b000000011101000010010110;
         rom[1101] = 24'b000000101010110011111101;
         rom[1102] = 24'b000000100101101100110010;
         rom[1103] = 24'b000000101000110010011111;
         rom[1104] = 24'b000000011000111110111000;
         rom[1105] = 24'b000000011010110000100101;
         rom[1106] = 24'b000000011011001101110101;
         rom[1107] = 24'b000000000111000101000010;
         rom[1108] = 24'b000000000101001111100010;
         rom[1109] = 24'b111111111110111100001110;
         rom[1110] = 24'b000000000001101110000110;
         rom[1111] = 24'b111111110011010010000111;
         rom[1112] = 24'b111111100100000111111101;
         rom[1113] = 24'b111111100011000010101100;
         rom[1114] = 24'b111111101001110111000101;
         rom[1115] = 24'b111111101001001100111111;
         rom[1116] = 24'b111111011000110000101101;
         rom[1117] = 24'b111111011011111101110001;
         rom[1118] = 24'b111111010110110110111101;
         rom[1119] = 24'b111111011111000000111011;
         rom[1120] = 24'b111111101001111110101000;
         rom[1121] = 24'b111111101001101000001101;
         rom[1122] = 24'b111111100110011000011011;
         rom[1123] = 24'b111111100000010111010110;
         rom[1124] = 24'b111111100110001000100011;
         rom[1125] = 24'b111111101101101001010001;
         rom[1126] = 24'b111111101101111101000110;
         rom[1127] = 24'b111111111011000101111110;
         rom[1128] = 24'b000000001011100110011000;
         rom[1129] = 24'b000000000000011001000110;
         rom[1130] = 24'b000000010101100010101100;
         rom[1131] = 24'b000000001111111000110011;
         rom[1132] = 24'b000000011000001010011101;
         rom[1133] = 24'b000000011010010010011101;
         rom[1134] = 24'b000000010101000001110001;
         rom[1135] = 24'b000000100110101010110110;
         rom[1136] = 24'b000000100001011101001001;
         rom[1137] = 24'b000000010110011101000110;
         rom[1138] = 24'b000000100110000011110001;
         rom[1139] = 24'b000000100110101011101010;
         rom[1140] = 24'b000000101110001011001110;
         rom[1141] = 24'b000000010100011001000011;
         rom[1142] = 24'b000000010000110110111100;
         rom[1143] = 24'b000000010000100110011100;
         rom[1144] = 24'b000000000110010011001110;
         rom[1145] = 24'b000000000100010000000100;
         rom[1146] = 24'b111111111111001101010100;
         rom[1147] = 24'b111111110111101011001100;
         rom[1148] = 24'b000000000001110100111000;
         rom[1149] = 24'b111111100010011111010111;
         rom[1150] = 24'b111111100101011111111001;
         rom[1151] = 24'b111111100011010100001100;
         rom[1152] = 24'b111111011000110011001011;
         rom[1153] = 24'b111111101101100010111001;
         rom[1154] = 24'b111111011001100100001100;
         rom[1155] = 24'b111111010110000010011010;
         rom[1156] = 24'b111111001111111001001110;
         rom[1157] = 24'b111111100010001101110110;
         rom[1158] = 24'b111111100011101010001000;
         rom[1159] = 24'b111111100010010001110100;
         rom[1160] = 24'b111111110001110000110111;
         rom[1161] = 24'b111111111000101101100001;
         rom[1162] = 24'b111111111001110110111101;
         rom[1163] = 24'b111111110101111110001001;
         rom[1164] = 24'b111111111110111000001110;
         rom[1165] = 24'b000000000101110100011001;
         rom[1166] = 24'b000000011000111101010110;
         rom[1167] = 24'b000000011110010110010001;
         rom[1168] = 24'b000000100010101001001101;
         rom[1169] = 24'b000000101001011000000011;
         rom[1170] = 24'b000000011000111001010110;
         rom[1171] = 24'b000000100010111001000000;
         rom[1172] = 24'b000000011000011000100110;
         rom[1173] = 24'b000000101111110010111010;
         rom[1174] = 24'b000000100010010001000101;
         rom[1175] = 24'b000000100010100110010001;
         rom[1176] = 24'b000000100101000001110000;
         rom[1177] = 24'b000000010110000011100101;
         rom[1178] = 24'b000000010101011110110100;
         rom[1179] = 24'b000000010001011000100010;
         rom[1180] = 24'b000000001100110011000101;
         rom[1181] = 24'b000000000100011100110110;
         rom[1182] = 24'b000000000000110101010110;
         rom[1183] = 24'b111111111000001000100110;
         rom[1184] = 24'b111111110011011010011001;
         rom[1185] = 24'b111111110001110001101110;
         rom[1186] = 24'b111111100110110101111010;
         rom[1187] = 24'b111111011010111000001010;
         rom[1188] = 24'b111111100001010011010000;
         rom[1189] = 24'b111111011110001101001111;
         rom[1190] = 24'b111111010011011100011010;
         rom[1191] = 24'b111111011000011110011110;
         rom[1192] = 24'b111111100011000101100101;
         rom[1193] = 24'b111111010111100011110011;
         rom[1194] = 24'b111111011110111101001001;
         rom[1195] = 24'b111111100000010000010111;
         rom[1196] = 24'b111111011111001000011111;
         rom[1197] = 24'b111111100011110111111111;
         rom[1198] = 24'b111111110011010011101000;
         rom[1199] = 24'b111111111000010000101111;
         rom[1200] = 24'b111111111101101010010011;
         rom[1201] = 24'b000000001110111011110001;
         rom[1202] = 24'b000000010010000011001101;
         rom[1203] = 24'b000000011100001110100010;
         rom[1204] = 24'b000000011111011000011000;
         rom[1205] = 24'b000000100011010001000110;
         rom[1206] = 24'b000000011100011000011100;
         rom[1207] = 24'b000000100000110000000110;
         rom[1208] = 24'b000000011010001011101101;
         rom[1209] = 24'b000000100101101111100101;
         rom[1210] = 24'b000000011110011000000011;
         rom[1211] = 24'b000000100100110111010110;
         rom[1212] = 24'b000000100000111110101111;
         rom[1213] = 24'b000000101100100000010110;
         rom[1214] = 24'b000000011111111010000011;
         rom[1215] = 24'b000000010000111010110100;
         rom[1216] = 24'b000000000100010100010000;
         rom[1217] = 24'b111111111010011011100000;
         rom[1218] = 24'b000000000011010110111011;
         rom[1219] = 24'b000000000011001001111000;
         rom[1220] = 24'b111111110100100101101111;
         rom[1221] = 24'b111111100111100111110110;
         rom[1222] = 24'b111111011100111010110111;
         rom[1223] = 24'b111111011100111111101010;
         rom[1224] = 24'b111111100011000111011101;
         rom[1225] = 24'b111111011100110011011011;
         rom[1226] = 24'b111111011010010110111110;
         rom[1227] = 24'b111111101010100110000001;
         rom[1228] = 24'b111111100010100100011100;
         rom[1229] = 24'b111111100011010100000000;
         rom[1230] = 24'b111111011011000010110000;
         rom[1231] = 24'b111111101111000100011110;
         rom[1232] = 24'b111111110100101111100011;
         rom[1233] = 24'b111111101101000001000110;
         rom[1234] = 24'b111111110100100111101111;
         rom[1235] = 24'b111111110010010100100100;
         rom[1236] = 24'b111111111101001100001001;
         rom[1237] = 24'b000000001010000011010101;
         rom[1238] = 24'b000000001010001110000000;
         rom[1239] = 24'b000000010000111010110100;
         rom[1240] = 24'b000000100001001001110100;
         rom[1241] = 24'b000000010100111001111001;
         rom[1242] = 24'b000000011000111100011101;
         rom[1243] = 24'b000000101101010001110110;
         rom[1244] = 24'b000000100011101100111101;
         rom[1245] = 24'b000000100010010010001001;
         rom[1246] = 24'b000000011101110101101111;
         rom[1247] = 24'b000000101011110011100111;
         rom[1248] = 24'b000000100011110001111000;
         rom[1249] = 24'b000000011110011110011111;
         rom[1250] = 24'b000000010110100001101101;
         rom[1251] = 24'b000000001111010011000011;
         rom[1252] = 24'b000000001010100110011100;
         rom[1253] = 24'b000000001011110010010001;
         rom[1254] = 24'b000000000111000000001100;
         rom[1255] = 24'b111111110110011011000101;
         rom[1256] = 24'b111111110111011100011110;
         rom[1257] = 24'b111111100101010000000111;
         rom[1258] = 24'b111111100111000100110011;
         rom[1259] = 24'b111111100011000001110001;
         rom[1260] = 24'b111111011001011011110001;
         rom[1261] = 24'b111111100000011011000110;
         rom[1262] = 24'b111111010111010100111010;
         rom[1263] = 24'b111111010110110001010110;
         rom[1264] = 24'b111111010111111001010011;
         rom[1265] = 24'b111111011011100100011000;
         rom[1266] = 24'b111111011010011101110010;
         rom[1267] = 24'b111111100010111101110100;
         rom[1268] = 24'b111111011100000100110100;
         rom[1269] = 24'b111111111000111010110011;
         rom[1270] = 24'b111111110100100101101001;
         rom[1271] = 24'b111111101000101100100101;
         rom[1272] = 24'b111111111001010100100100;
         rom[1273] = 24'b111111111111111001110011;
         rom[1274] = 24'b000000010001100010101101;
         rom[1275] = 24'b000000001111010110010010;
         rom[1276] = 24'b000000011000101110101010;
         rom[1277] = 24'b000000010011010110100110;
         rom[1278] = 24'b000000011101110110100001;
         rom[1279] = 24'b000000011111101111110100;
         rom[1280] = 24'b000000100010001100110111;
         rom[1281] = 24'b000000101001011101000000;
         rom[1282] = 24'b000000011011000101100101;
         rom[1283] = 24'b000000100011100101111000;
         rom[1284] = 24'b000000110100101101110000;
         rom[1285] = 24'b000000011100111111010101;
         rom[1286] = 24'b000000100101110100100101;
         rom[1287] = 24'b000000010111011000011110;
         rom[1288] = 24'b000000001000101100100101;
         rom[1289] = 24'b000000001000010101001010;
         rom[1290] = 24'b000000000111000101010011;
         rom[1291] = 24'b111111111010000110100111;
         rom[1292] = 24'b111111111011010001101010;
         rom[1293] = 24'b111111111011111100100010;
         rom[1294] = 24'b111111110011011000001100;
         rom[1295] = 24'b111111011111001000010000;
         rom[1296] = 24'b111111101000000001100100;
         rom[1297] = 24'b111111101100010011011001;
         rom[1298] = 24'b111111100010110010101001;
         rom[1299] = 24'b111111011110110001011000;
         rom[1300] = 24'b111111001111010010011111;
         rom[1301] = 24'b111111011101000001110110;
         rom[1302] = 24'b111111110001001101010001;
         rom[1303] = 24'b111111111001110000000110;
         rom[1304] = 24'b111111111111011011100111;
         rom[1305] = 24'b000000001110010101101001;
         rom[1306] = 24'b000000010011111110110100;
         rom[1307] = 24'b000000101000100111101111;
         rom[1308] = 24'b000000101000111011011001;
         rom[1309] = 24'b000001000100110010001101;
         rom[1310] = 24'b000001010010000000001110;
         rom[1311] = 24'b000001011001100110001111;
         rom[1312] = 24'b000001110000101100100101;
         rom[1313] = 24'b000001101110001001101100;
         rom[1314] = 24'b000010000100001001011100;
         rom[1315] = 24'b000010001111110011011111;
         rom[1316] = 24'b000010011011101000001000;
         rom[1317] = 24'b000010101010010011001110;
         rom[1318] = 24'b000010101100110010110010;
         rom[1319] = 24'b000010110100001011011110;
         rom[1320] = 24'b000010110111000001000000;
         rom[1321] = 24'b000010110010000100000001;
         rom[1322] = 24'b000010111110001110001100;
         rom[1323] = 24'b000010111011111000111111;
         rom[1324] = 24'b000011000010111100011111;
         rom[1325] = 24'b000011001001100010101100;
         rom[1326] = 24'b000010111111111010110011;
         rom[1327] = 24'b000011000100110111011001;
         rom[1328] = 24'b000010111101110111111101;
         rom[1329] = 24'b000011010010001100000101;
         rom[1330] = 24'b000011010010000110001010;
         rom[1331] = 24'b000011001100001100110101;
         rom[1332] = 24'b000011001010100000101000;
         rom[1333] = 24'b000011001101001101011010;
         rom[1334] = 24'b000011010111001000101000;
         rom[1335] = 24'b000011011001011011100101;
         rom[1336] = 24'b000011010001010110010100;
         rom[1337] = 24'b000011110010010110010001;
         rom[1338] = 24'b000011110001000110001110;
         rom[1339] = 24'b000011110101011011000011;
         rom[1340] = 24'b000100001100011010101111;
         rom[1341] = 24'b000100010000111001010101;
         rom[1342] = 24'b000100010011100011100011;
         rom[1343] = 24'b000100100111010010010000;
         rom[1344] = 24'b000100111001001001011100;
         rom[1345] = 24'b000100111111110100111011;
         rom[1346] = 24'b000101011011111111010100;
         rom[1347] = 24'b000101100001100001110101;
         rom[1348] = 24'b000101101011100101110010;
         rom[1349] = 24'b000101111000101110010100;
         rom[1350] = 24'b000110010011011001001000;
         rom[1351] = 24'b000110000110011001111110;
         rom[1352] = 24'b000110011111000110110000;
         rom[1353] = 24'b000110110110110110011011;
         rom[1354] = 24'b000110100110000111110011;
         rom[1355] = 24'b000110111001001111000011;
         rom[1356] = 24'b000110110110010110000011;
         rom[1357] = 24'b000110111111000110101100;
         rom[1358] = 24'b000111000010010111001111;
         rom[1359] = 24'b000111000001101101101110;
         rom[1360] = 24'b000111000011110001010101;
         rom[1361] = 24'b000111010100110110001000;
         rom[1362] = 24'b000111010101100000111100;
         rom[1363] = 24'b000111010010010010011110;
         rom[1364] = 24'b000111010000110101110101;
         rom[1365] = 24'b000111001101001000100111;
         rom[1366] = 24'b000111001010000001011011;
         rom[1367] = 24'b000111001100100000111000;
         rom[1368] = 24'b000111100110100001010000;
         rom[1369] = 24'b000111011000110110110000;
         rom[1370] = 24'b000111100001101010111011;
         rom[1371] = 24'b000111100000110101001011;
         rom[1372] = 24'b000111100100101100010101;
         rom[1373] = 24'b000111111001100000110011;
         rom[1374] = 24'b000111110011111011011111;
         rom[1375] = 24'b001000010000011000001110;
         rom[1376] = 24'b001000000110001110000000;
         rom[1377] = 24'b001000000111101101100001;
         rom[1378] = 24'b001000011101100001100001;
         rom[1379] = 24'b001000100111100101110110;
         rom[1380] = 24'b001001000010101011111101;
         rom[1381] = 24'b001001001011101110010111;
         rom[1382] = 24'b001001010001000010110100;
         rom[1383] = 24'b001001100100011100111010;
         rom[1384] = 24'b001001110011110100000111;
         rom[1385] = 24'b001001111100101010000110;
         rom[1386] = 24'b001010010000001111100111;
         rom[1387] = 24'b001010011001001100100001;
         rom[1388] = 24'b001010011101101011010001;
         rom[1389] = 24'b001010010011010100111110;
         rom[1390] = 24'b001010010101011000100111;
         rom[1391] = 24'b001001111110111100010010;
         rom[1392] = 24'b001001111111101100100001;
         rom[1393] = 24'b001001110000011011110101;
         rom[1394] = 24'b001001101010001111011101;
         rom[1395] = 24'b001001101011000011011101;
         rom[1396] = 24'b001001011001000001110110;
         rom[1397] = 24'b001001010010011001001111;
         rom[1398] = 24'b001001000000011010011001;
         rom[1399] = 24'b001000101011001010000000;
         rom[1400] = 24'b001000100010100001010011;
         rom[1401] = 24'b001000001010010010011001;
         rom[1402] = 24'b000111111011101001001000;
         rom[1403] = 24'b001000001100010110000101;
         rom[1404] = 24'b000111101000111001111010;
         rom[1405] = 24'b000111100100101001001111;
         rom[1406] = 24'b000111001110110000110101;
         rom[1407] = 24'b000111010100011111001001;
         rom[1408] = 24'b000111001001011111001110;
         rom[1409] = 24'b000111000011010100100000;
         rom[1410] = 24'b000110110111010100100111;
         rom[1411] = 24'b000110101000011001111001;
         rom[1412] = 24'b000110111011101010001000;
         rom[1413] = 24'b000110011010100111001111;
         rom[1414] = 24'b000110011111011110010101;
         rom[1415] = 24'b000110101001011010100010;
         rom[1416] = 24'b000110011111110101111000;
         rom[1417] = 24'b000110100110000101100010;
         rom[1418] = 24'b000110100100110110111011;
         rom[1419] = 24'b000110011000100110001000;
         rom[1420] = 24'b000110100100001001111110;
         rom[1421] = 24'b000110011001110100101101;
         rom[1422] = 24'b000110010010000011010110;
         rom[1423] = 24'b000110011110001110101010;
         rom[1424] = 24'b000110011011111100111110;
         rom[1425] = 24'b000110010011111100010010;
         rom[1426] = 24'b000110001001110001110000;
         rom[1427] = 24'b000101111010010100100010;
         rom[1428] = 24'b000110000000000110001101;
         rom[1429] = 24'b000101110110101000100101;
         rom[1430] = 24'b000101100111111101001000;
         rom[1431] = 24'b000101011101101100100111;
         rom[1432] = 24'b000101010111010011110000;
         rom[1433] = 24'b000101000100100100100010;
         rom[1434] = 24'b000100111101101011111101;
         rom[1435] = 24'b000100101101101011110011;
         rom[1436] = 24'b000100100010011011101001;
         rom[1437] = 24'b000100010011011001011100;
         rom[1438] = 24'b000100000111100010010110;
         rom[1439] = 24'b000011111010000011011111;
         rom[1440] = 24'b000011110011011000111110;
         rom[1441] = 24'b000011101010001110100100;
         rom[1442] = 24'b000011011010110000101111;
         rom[1443] = 24'b000011000100001101010111;
         rom[1444] = 24'b000010111101101100001001;
         rom[1445] = 24'b000010110001011000111101;
         rom[1446] = 24'b000010110101101111011111;
         rom[1447] = 24'b000010101010010011110000;
         rom[1448] = 24'b000010101101100000011111;
         rom[1449] = 24'b000010011001110110000111;
         rom[1450] = 24'b000010100011100100011101;
         rom[1451] = 24'b000010011110111011101010;
         rom[1452] = 24'b000010001100001100001000;
         rom[1453] = 24'b000010100110001001101101;
         rom[1454] = 24'b000010011010110110001001;
         rom[1455] = 24'b000010011001101011010101;
         rom[1456] = 24'b000010010100111010101001;
         rom[1457] = 24'b000010010101000100101010;
         rom[1458] = 24'b000010010010101000011000;
         rom[1459] = 24'b000010000110110000000000;
         rom[1460] = 24'b000010000011011000101101;
         rom[1461] = 24'b000010000011100110101000;
         rom[1462] = 24'b000010010101000011110011;
         rom[1463] = 24'b000010000010001011010110;
         rom[1464] = 24'b000001111011111010010111;
         rom[1465] = 24'b000001101100011011100101;
         rom[1466] = 24'b000001101011111010011001;
         rom[1467] = 24'b000001011110110111100001;
         rom[1468] = 24'b000001000111011100010111;
         rom[1469] = 24'b000001000111100001000101;
         rom[1470] = 24'b000000111100000011000111;
         rom[1471] = 24'b000000011110011010111001;
         rom[1472] = 24'b000000011110110000010110;
         rom[1473] = 24'b000000000001011011100110;
         rom[1474] = 24'b111111111100101101011000;
         rom[1475] = 24'b111111101100010001110011;
         rom[1476] = 24'b111111100110110001100001;
         rom[1477] = 24'b111111100010000001010110;
         rom[1478] = 24'b111111010100101101010100;
         rom[1479] = 24'b111111001011000111111110;
         rom[1480] = 24'b111110110110011011111000;
         rom[1481] = 24'b111110101011101100011011;
         rom[1482] = 24'b111110110100010001011101;
         rom[1483] = 24'b111110100111000110100110;
         rom[1484] = 24'b111110011110000010001000;
         rom[1485] = 24'b111110011101010101111001;
         rom[1486] = 24'b111110000110101100000101;
         rom[1487] = 24'b111110010011001010100111;
         rom[1488] = 24'b111110011000111000111011;
         rom[1489] = 24'b111110101001011001100010;
         rom[1490] = 24'b111110101011110000111000;
         rom[1491] = 24'b111110111011110100100000;
         rom[1492] = 24'b111111010100100111001011;
         rom[1493] = 24'b111111011011010000111111;
         rom[1494] = 24'b111111100011000110111010;
         rom[1495] = 24'b111111110111011000000010;
         rom[1496] = 24'b111111110001110001011001;
         rom[1497] = 24'b000000001000101101000001;
         rom[1498] = 24'b000000010011011000111011;
         rom[1499] = 24'b000000011010100101000000;
         rom[1500] = 24'b000000100010101100111010;
         rom[1501] = 24'b000000100010000110111111;
         rom[1502] = 24'b000000101001010000000111;
         rom[1503] = 24'b000000100011110101111111;
         rom[1504] = 24'b000000100001100110011000;
         rom[1505] = 24'b000000011010101010101101;
         rom[1506] = 24'b000000001010011011001011;
         rom[1507] = 24'b000000011000110101110011;
         rom[1508] = 24'b111111110111010010011100;
         rom[1509] = 24'b000000000111001110001101;
         rom[1510] = 24'b111111111100010001000101;
         rom[1511] = 24'b111111101101001111010001;
         rom[1512] = 24'b111111110000000010111010;
         rom[1513] = 24'b111111110000000010111011;
         rom[1514] = 24'b111111011110110000011011;
         rom[1515] = 24'b111111100100110110111111;
         rom[1516] = 24'b111111011100000011001111;
         rom[1517] = 24'b111111010110100110001100;
         rom[1518] = 24'b111111011111100101100111;
         rom[1519] = 24'b111111011110111111010011;
         rom[1520] = 24'b111111011110000100100100;
         rom[1521] = 24'b111111100110010100010111;
         rom[1522] = 24'b111111101011010010100111;
         rom[1523] = 24'b111111100110110011110101;
         rom[1524] = 24'b111111100111101000011111;
         rom[1525] = 24'b111111110100110011001011;
         rom[1526] = 24'b111111110100110101011100;
         rom[1527] = 24'b111111111000111010111001;
         rom[1528] = 24'b000000000110000000011101;
         rom[1529] = 24'b000000000011000100010110;
         rom[1530] = 24'b000000011111001110010010;
         rom[1531] = 24'b000000011111100101111001;
         rom[1532] = 24'b000000011100000111001101;
         rom[1533] = 24'b000000011110110100100110;
         rom[1534] = 24'b000000100000000111010011;
         rom[1535] = 24'b000000101011110111001001;
         rom[1536] = 24'b000000100101010100100001;
         rom[1537] = 24'b000000011111001110001000;
         rom[1538] = 24'b000000100000011101100001;
         rom[1539] = 24'b000000100101111111100000;
         rom[1540] = 24'b000000100101010101101111;
         rom[1541] = 24'b000000011000100010100100;
         rom[1542] = 24'b000000010001101111110111;
         rom[1543] = 24'b000000001101010001001110;
         rom[1544] = 24'b000000010010001111011110;
         rom[1545] = 24'b111111110100111100011011;
         rom[1546] = 24'b111111111100101000011110;
         rom[1547] = 24'b111111111100001000010011;
         rom[1548] = 24'b111111100001001011001110;
         rom[1549] = 24'b111111101110100101001110;
         rom[1550] = 24'b111111101100001110111110;
         rom[1551] = 24'b111111010000101100110001;
         rom[1552] = 24'b111111011001100111010111;
         rom[1553] = 24'b111111010111010101110111;
         rom[1554] = 24'b111111001111010101100101;
         rom[1555] = 24'b111111011011011111000110;
         rom[1556] = 24'b111111100001010011110111;
         rom[1557] = 24'b111111101000000011100000;
         rom[1558] = 24'b111111110100001101001011;
         rom[1559] = 24'b111111110010101010000111;
         rom[1560] = 24'b111111100101011011101001;
         rom[1561] = 24'b111111101010110101000001;
         rom[1562] = 24'b111111111001100100011110;
         rom[1563] = 24'b111111111100100000000000;
         rom[1564] = 24'b000000001000101101101001;
         rom[1565] = 24'b000000000110010001111010;
         rom[1566] = 24'b000000001010000001000000;
         rom[1567] = 24'b000000010110011100110101;
         rom[1568] = 24'b000000001101010111101100;
         rom[1569] = 24'b000000011100111110011010;
         rom[1570] = 24'b000000100110110101010001;
         rom[1571] = 24'b000000101010101111010010;
         rom[1572] = 24'b000000100000000000100010;
         rom[1573] = 24'b000000100111110110100110;
         rom[1574] = 24'b000000100111001111111011;
         rom[1575] = 24'b000000100010001011111001;
         rom[1576] = 24'b000000011000000110010110;
         rom[1577] = 24'b000000010000111100010101;
         rom[1578] = 24'b000000001101000100110100;
         rom[1579] = 24'b000000010100101010101101;
         rom[1580] = 24'b000000010011101010110001;
         rom[1581] = 24'b000000001011001100010100;
         rom[1582] = 24'b000000000001100100110001;
         rom[1583] = 24'b111111110000101101011011;
         rom[1584] = 24'b111111101111101000110100;
         rom[1585] = 24'b111111101100001000111011;
         rom[1586] = 24'b111111011110010101001100;
         rom[1587] = 24'b111111100101111000101100;
         rom[1588] = 24'b111111100111110011110101;
         rom[1589] = 24'b111111010010000111000011;
         rom[1590] = 24'b111111011011000000100111;
         rom[1591] = 24'b111111011111000111000111;
         rom[1592] = 24'b111111011000100011000000;
         rom[1593] = 24'b111111011100000000101111;
         rom[1594] = 24'b111111101011010110111001;
         rom[1595] = 24'b111111100011000001010011;
         rom[1596] = 24'b111111101000101101000010;
         rom[1597] = 24'b000000000010011111101110;
         rom[1598] = 24'b111111101001100010110000;
         rom[1599] = 24'b111111110100010000010011;
         rom[1600] = 24'b111111110110111000011101;
         rom[1601] = 24'b000000000100010110001100;
         rom[1602] = 24'b000000010110000000100100;
         rom[1603] = 24'b000000010000100110011010;
         rom[1604] = 24'b000000010110110111010111;
         rom[1605] = 24'b000000100000010100011011;
         rom[1606] = 24'b000000011101110011111011;
         rom[1607] = 24'b000000101010011101011111;
         rom[1608] = 24'b000000100110100000110010;
         rom[1609] = 24'b000000100010110101011110;
         rom[1610] = 24'b000000011100001011000000;
         rom[1611] = 24'b000000011111100111010111;
         rom[1612] = 24'b000000010101111101110110;
         rom[1613] = 24'b000000010101011101011011;
         rom[1614] = 24'b000000001100110010101011;
         rom[1615] = 24'b000000010001110001101010;
         rom[1616] = 24'b000000001100100000100011;
         rom[1617] = 24'b000000000010110101101100;
         rom[1618] = 24'b111111111011110000010101;
         rom[1619] = 24'b111111111111111000011101;
         rom[1620] = 24'b111111110011001111100101;
         rom[1621] = 24'b111111111001001101110111;
         rom[1622] = 24'b111111101010100111000000;
         rom[1623] = 24'b111111110001110111100000;
         rom[1624] = 24'b111111100101001001111001;
         rom[1625] = 24'b111111100010110111000001;
         rom[1626] = 24'b111111011111001110001001;
         rom[1627] = 24'b111111101000010100010011;
         rom[1628] = 24'b111111101000010000010111;
         rom[1629] = 24'b111111011110111001100001;
         rom[1630] = 24'b111111011110011001100000;
         rom[1631] = 24'b111111011111011010010111;
         rom[1632] = 24'b111111110010011011010011;
         rom[1633] = 24'b111111111000111100111111;
         rom[1634] = 24'b111111101100011111011110;
         rom[1635] = 24'b111111100101000110100000;
         rom[1636] = 24'b111111110101010101101110;
         rom[1637] = 24'b000000001111111100000101;
         rom[1638] = 24'b000000000110011001111101;
         rom[1639] = 24'b000000010001111001111001;
         rom[1640] = 24'b000000010011101100110110;
         rom[1641] = 24'b000000100101110111100111;
         rom[1642] = 24'b000000101111110101010000;
         rom[1643] = 24'b000000100111110111000100;
         rom[1644] = 24'b000000111010111101011001;
         rom[1645] = 24'b000001001001000100001010;
         rom[1646] = 24'b000001000011010101010101;
         rom[1647] = 24'b000001000011100000000001;
         rom[1648] = 24'b000000110010010000001010;
         rom[1649] = 24'b000001000011001011000010;
         rom[1650] = 24'b000001000100010100001001;
         rom[1651] = 24'b000001000101101001000110;
         rom[1652] = 24'b000000111111010001011100;
         rom[1653] = 24'b000000110100111110011011;
         rom[1654] = 24'b000000111000100101000101;
         rom[1655] = 24'b000000101001011100110011;
         rom[1656] = 24'b000000101010101100111010;
         rom[1657] = 24'b000000011100101000101001;
         rom[1658] = 24'b000000011001000000110010;
         rom[1659] = 24'b000000100001001001010110;
         rom[1660] = 24'b000000010011000100000101;
         rom[1661] = 24'b000000011100010011000001;
         rom[1662] = 24'b000000001110101001101000;
         rom[1663] = 24'b000000010010001110010101;
         rom[1664] = 24'b000000011010011011011000;
         rom[1665] = 24'b000000001001110011111000;
         rom[1666] = 24'b000000011000000110110001;
         rom[1667] = 24'b000000101100101010101100;
         rom[1668] = 24'b000000011100100010111100;
         rom[1669] = 24'b000000111111001101000001;
         rom[1670] = 24'b000000101111110111111110;
         rom[1671] = 24'b000000110110100001001110;
         rom[1672] = 24'b000000111010100010100001;
         rom[1673] = 24'b000000111111101101010101;
         rom[1674] = 24'b000001001110110100101010;
         rom[1675] = 24'b000001010101011010110110;
         rom[1676] = 24'b000001100011101100011001;
         rom[1677] = 24'b000001011111110001001001;
         rom[1678] = 24'b000001100111001110011010;
         rom[1679] = 24'b000001100010101001011110;
         rom[1680] = 24'b000001101111111100010010;
         rom[1681] = 24'b000001111110000000011010;
         rom[1682] = 24'b000001101110011100011111;
         rom[1683] = 24'b000001100010000001111111;
         rom[1684] = 24'b000001101101100100110100;
         rom[1685] = 24'b000001011101000100010011;
         rom[1686] = 24'b000001100001110001011111;
         rom[1687] = 24'b000001110000000000111010;
         rom[1688] = 24'b000001011001100000011111;
         rom[1689] = 24'b000001100010010101001101;
         rom[1690] = 24'b000001011110000101000111;
         rom[1691] = 24'b000001011011011011100010;
         rom[1692] = 24'b000001010000111100011001;
         rom[1693] = 24'b000001000001101011100111;
         rom[1694] = 24'b000001001000111010110011;
         rom[1695] = 24'b000001000011011010011001;
         rom[1696] = 24'b000000111110101110001011;
         rom[1697] = 24'b000000111011101111001011;
         rom[1698] = 24'b000000110011111000111101;
         rom[1699] = 24'b000000111100011000111000;
         rom[1700] = 24'b000000110101001010010111;
         rom[1701] = 24'b000001000010100100011111;
         rom[1702] = 24'b000000111010111111111011;
         rom[1703] = 24'b000000111011001011110001;
         rom[1704] = 24'b000001001000101101110101;
         rom[1705] = 24'b000000111111001111010111;
         rom[1706] = 24'b000001001101111100000011;
         rom[1707] = 24'b000001010011100111111101;
         rom[1708] = 24'b000001010101010110110011;
         rom[1709] = 24'b000001101011010110110011;
         rom[1710] = 24'b000001101110110010010000;
         rom[1711] = 24'b000001110110010000000111;
         rom[1712] = 24'b000001101100001000111000;
         rom[1713] = 24'b000001111111100011010000;
         rom[1714] = 24'b000010000101000001010000;
         rom[1715] = 24'b000010010011101001010111;
         rom[1716] = 24'b000010001000011010101100;
         rom[1717] = 24'b000010000010110100111101;
         rom[1718] = 24'b000010000010001011000011;
         rom[1719] = 24'b000010000111001110101110;
         rom[1720] = 24'b000010000111100010101010;
         rom[1721] = 24'b000010000111100011111100;
         rom[1722] = 24'b000010000110110111100011;
         rom[1723] = 24'b000001111011111011000000;
         rom[1724] = 24'b000001110110100011101100;
         rom[1725] = 24'b000001110100001011011010;
         rom[1726] = 24'b000001100110111110110111;
         rom[1727] = 24'b000001100000011010001111;
         rom[1728] = 24'b000001101110011000011011;
         rom[1729] = 24'b000001011110100111001100;
         rom[1730] = 24'b000001100010101111111111;
         rom[1731] = 24'b000001010010011000011111;
         rom[1732] = 24'b000001010001000111111001;
         rom[1733] = 24'b000001001101101011110000;
         rom[1734] = 24'b000001000100101100010100;
         rom[1735] = 24'b000001010101011100000010;
         rom[1736] = 24'b000001000100011111010110;
         rom[1737] = 24'b000001000001010110000101;
         rom[1738] = 24'b000001000011000111100011;
         rom[1739] = 24'b000001000110010000101100;
         rom[1740] = 24'b000001000111101101010101;
         rom[1741] = 24'b000001011011110100100101;
         rom[1742] = 24'b000001011000011111110100;
         rom[1743] = 24'b000001110001010010011111;
         rom[1744] = 24'b000001100100011101001011;
         rom[1745] = 24'b000001111000001100101100;
         rom[1746] = 24'b000001101101001100010100;
         rom[1747] = 24'b000001111011011011101100;
         rom[1748] = 24'b000001111001110001000000;
         rom[1749] = 24'b000001111111100111101010;
         rom[1750] = 24'b000010000100110100010111;
         rom[1751] = 24'b000010001110010111101110;
         rom[1752] = 24'b000010010111110001011000;
         rom[1753] = 24'b000010010010001101010110;
         rom[1754] = 24'b000010000110001000010111;
         rom[1755] = 24'b000010001001010100010011;
         rom[1756] = 24'b000010010100111010001010;
         rom[1757] = 24'b000010000111100011100100;
         rom[1758] = 24'b000010011000011010110111;
         rom[1759] = 24'b000010011100011011000010;
         rom[1760] = 24'b000010000001011100111100;
         rom[1761] = 24'b000010010001001010100110;
         rom[1762] = 24'b000001111111001111101000;
         rom[1763] = 24'b000001101111001001110111;
         rom[1764] = 24'b000001100110010100001111;
         rom[1765] = 24'b000001101110001100000000;
         rom[1766] = 24'b000001011100000011101000;
         rom[1767] = 24'b000001011011111101011111;
         rom[1768] = 24'b000001011110110000000111;
         rom[1769] = 24'b000001011000011011011110;
         rom[1770] = 24'b000001010100111000001011;
         rom[1771] = 24'b000001011010110110011100;
         rom[1772] = 24'b000001010111101100000010;
         rom[1773] = 24'b000001000111000001101101;
         rom[1774] = 24'b000001011100001001011010;
         rom[1775] = 24'b000001010110000101111101;
         rom[1776] = 24'b000001011000111100000001;
         rom[1777] = 24'b000001100001101010110110;
         rom[1778] = 24'b000001011011001010100110;
         rom[1779] = 24'b000001100000000110011101;
         rom[1780] = 24'b000001111010101110101001;
         rom[1781] = 24'b000001110101010110101010;
         rom[1782] = 24'b000001110011100001100000;
         rom[1783] = 24'b000001110101011001011101;
         rom[1784] = 24'b000010010101111110011111;
         rom[1785] = 24'b000010001000110110010000;
         rom[1786] = 24'b000010001110010000111101;
         rom[1787] = 24'b000010001000001110011101;
         rom[1788] = 24'b000010010001100001010011;
         rom[1789] = 24'b000010010110111011001010;
         rom[1790] = 24'b000010101000011001001111;
         rom[1791] = 24'b000010011001101000000000;
         rom[1792] = 24'b000010011101101100000110;
         rom[1793] = 24'b000010011001111010100101;
         rom[1794] = 24'b000010010010001101000100;
         rom[1795] = 24'b000010010011101111111111;
         rom[1796] = 24'b000010001010111011000111;
         rom[1797] = 24'b000010010001001101011111;
         rom[1798] = 24'b000001111100110000110010;
         rom[1799] = 24'b000001110111011100001010;
         rom[1800] = 24'b000001110101001001110111;
         rom[1801] = 24'b000001110000100001010000;
         rom[1802] = 24'b000001100111001010010001;
         rom[1803] = 24'b000001100111010110001111;
         rom[1804] = 24'b000001100010001111111101;
         rom[1805] = 24'b000001010111111100000001;
         rom[1806] = 24'b000001010001111001111010;
         rom[1807] = 24'b000001100101000101101101;
         rom[1808] = 24'b000001011111010010001101;
         rom[1809] = 24'b000001010111010110100010;
         rom[1810] = 24'b000001001101100101110000;
         rom[1811] = 24'b000001011000010001100101;
         rom[1812] = 24'b000001100110000001001000;
         rom[1813] = 24'b000001010001001000011111;
         rom[1814] = 24'b000001011001101111101010;
         rom[1815] = 24'b000001100011111000010011;
         rom[1816] = 24'b000001110010010011001101;
         rom[1817] = 24'b000001110010000111010000;
         rom[1818] = 24'b000001101100100101011100;
         rom[1819] = 24'b000010000111100111101101;
         rom[1820] = 24'b000001110001001010101001;
         rom[1821] = 24'b000010010010010001000111;
         rom[1822] = 24'b000010011011100010001111;
         rom[1823] = 24'b000010011010100001110001;
         rom[1824] = 24'b000010010010011101101111;
         rom[1825] = 24'b000010011111001110111100;
         rom[1826] = 24'b000010100100011111110001;
         rom[1827] = 24'b000010010000111100010001;
         rom[1828] = 24'b000010001100111111000000;
         rom[1829] = 24'b000010100101101010100011;
         rom[1830] = 24'b000010001111101100000010;
         rom[1831] = 24'b000010010111101011001111;
         rom[1832] = 24'b000010001110010111101000;
         rom[1833] = 24'b000010001101101101111110;
         rom[1834] = 24'b000001111101011111110100;
         rom[1835] = 24'b000001111110100111111001;
         rom[1836] = 24'b000001111100001010010000;
         rom[1837] = 24'b000001110100000010111110;
         rom[1838] = 24'b000001110101011111010110;
         rom[1839] = 24'b000001110110100000101010;
         rom[1840] = 24'b000001100000011010000100;
         rom[1841] = 24'b000001100000101010001001;
         rom[1842] = 24'b000001011010010101111010;
         rom[1843] = 24'b000001010101001110101110;
         rom[1844] = 24'b000001011001011111100011;
         rom[1845] = 24'b000001001010000010011111;
         rom[1846] = 24'b000001100000010010110110;
         rom[1847] = 24'b000001011000000000010110;
         rom[1848] = 24'b000001001000111010100000;
         rom[1849] = 24'b000001011001000001011100;
         rom[1850] = 24'b000001100001001001100110;
         rom[1851] = 24'b000001011011001000110100;
         rom[1852] = 24'b000001111000011010011001;
         rom[1853] = 24'b000001101000001111001101;
         rom[1854] = 24'b000001101010001010100000;
         rom[1855] = 24'b000001111110110001110000;
         rom[1856] = 24'b000001111011001100000000;
         rom[1857] = 24'b000010000110111011100110;
         rom[1858] = 24'b000010001101001100101010;
         rom[1859] = 24'b000010010111001100010000;
         rom[1860] = 24'b000010010001110001000100;
         rom[1861] = 24'b000010011101101010111111;
         rom[1862] = 24'b000010010011111101100100;
         rom[1863] = 24'b000010010100000011001110;
         rom[1864] = 24'b000010011111001101000111;
         rom[1865] = 24'b000010011001100100010101;
         rom[1866] = 24'b000010001111100111111101;
         rom[1867] = 24'b000010011001000000110111;
         rom[1868] = 24'b000010011001111111001011;
         rom[1869] = 24'b000010001101101000001000;
         rom[1870] = 24'b000010001000010110001001;
         rom[1871] = 24'b000001110101001000110101;
         rom[1872] = 24'b000010000000011000100000;
         rom[1873] = 24'b000001110110011000100111;
         rom[1874] = 24'b000001110011001100011100;
         rom[1875] = 24'b000001011010000100001010;
         rom[1876] = 24'b000001101101011011101100;
         rom[1877] = 24'b000001101011111110101000;
         rom[1878] = 24'b000001011001101111100100;
         rom[1879] = 24'b000001100011111011000010;
         rom[1880] = 24'b000001011000010111001011;
         rom[1881] = 24'b000001010100000111100010;
         rom[1882] = 24'b000001001000111100010001;
         rom[1883] = 24'b000001010100000100100010;
         rom[1884] = 24'b000001011100010100000011;
         rom[1885] = 24'b000001001110001110001011;
         rom[1886] = 24'b000001010100100110000000;
         rom[1887] = 24'b000001100100011010100101;
         rom[1888] = 24'b000001100011010011110100;
         rom[1889] = 24'b000001011110000001010110;
         rom[1890] = 24'b000001111010000010110000;
         rom[1891] = 24'b000001101001010111010011;
         rom[1892] = 24'b000001111000111110010100;
         rom[1893] = 24'b000001110001101110100010;
         rom[1894] = 24'b000010001000000101111010;
         rom[1895] = 24'b000010001110001000010000;
         rom[1896] = 24'b000010000001011000101111;
         rom[1897] = 24'b000010000000011000000101;
         rom[1898] = 24'b000010001001100110000001;
         rom[1899] = 24'b000010010010011010011100;
         rom[1900] = 24'b000010001110101001001000;
         rom[1901] = 24'b000010001011011111110110;
         rom[1902] = 24'b000010010110001100011000;
         rom[1903] = 24'b000010010001100001101111;
         rom[1904] = 24'b000001110111011001110010;
         rom[1905] = 24'b000010001011101101110101;
         rom[1906] = 24'b000010000001010100101110;
         rom[1907] = 24'b000010000100110001101101;
         rom[1908] = 24'b000001100111111101011011;
         rom[1909] = 24'b000001100111110111111111;
         rom[1910] = 24'b000001011101111000000101;
         rom[1911] = 24'b000001100001011101100111;
         rom[1912] = 24'b000001001111010111100110;
         rom[1913] = 24'b000001010111111101111100;
         rom[1914] = 24'b000001000110011111010011;
         rom[1915] = 24'b000001001011101101001011;
         rom[1916] = 24'b000001000001101111000101;
         rom[1917] = 24'b000000111100000101000011;
         rom[1918] = 24'b000000110010111111010111;
         rom[1919] = 24'b000000111110100100010110;
         rom[1920] = 24'b000001000000100001000111;
         rom[1921] = 24'b000001000111110010001101;
         rom[1922] = 24'b000000111010011011000000;
         rom[1923] = 24'b000001010000001100001011;
         rom[1924] = 24'b000001011001000011101100;
         rom[1925] = 24'b000001011101000010100000;
         rom[1926] = 24'b000001100000000111011010;
         rom[1927] = 24'b000001011110010100010011;
         rom[1928] = 24'b000001010100110110000101;
         rom[1929] = 24'b000001101100101101111000;
         rom[1930] = 24'b000001111000000100111000;
         rom[1931] = 24'b000001111000110011000001;
         rom[1932] = 24'b000001111011101000100110;
         rom[1933] = 24'b000001110101010010101101;
         rom[1934] = 24'b000010001000000001001100;
         rom[1935] = 24'b000010001101111001101101;
         rom[1936] = 24'b000010001101111011010101;
         rom[1937] = 24'b000001111101101011010101;
         rom[1938] = 24'b000010001000010111011100;
         rom[1939] = 24'b000001111001001100010110;
         rom[1940] = 24'b000001110110100101011010;
         rom[1941] = 24'b000001110000110001101010;
         rom[1942] = 24'b000001101000100111111011;
         rom[1943] = 24'b000001101110001011101111;
         rom[1944] = 24'b000001101111001110101011;
         rom[1945] = 24'b000001010011000010111100;
         rom[1946] = 24'b000001001000100101011001;
         rom[1947] = 24'b000001001011100111100100;
         rom[1948] = 24'b000001001001100000100011;
         rom[1949] = 24'b000000111101001011011101;
         rom[1950] = 24'b000000111001000011100001;
         rom[1951] = 24'b000001000110011010011101;
         rom[1952] = 24'b000000101111111011010001;
         rom[1953] = 24'b000000101010111101110011;
         rom[1954] = 24'b000000101100100000110110;
         rom[1955] = 24'b000000101010001001001110;
         rom[1956] = 24'b000000011111110000010100;
         rom[1957] = 24'b000000110010000100111010;
         rom[1958] = 24'b000000110100000111001101;
         rom[1959] = 24'b000001000010010110011000;
         rom[1960] = 24'b000000110000000011101101;
         rom[1961] = 24'b000000111101001110101101;
         rom[1962] = 24'b000000111110001000011000;
         rom[1963] = 24'b000001001011001001100101;
         rom[1964] = 24'b000001001111101000011101;
         rom[1965] = 24'b000000111011011011010011;
         rom[1966] = 24'b000001001101011110110000;
         rom[1967] = 24'b000001011100111101111111;
         rom[1968] = 24'b000001011110011000001010;
         rom[1969] = 24'b000001100010011010100011;
         rom[1970] = 24'b000001101000011101010010;
         rom[1971] = 24'b000001101110101101111010;
         rom[1972] = 24'b000001011010000000010001;
         rom[1973] = 24'b000001100101011001011100;
         rom[1974] = 24'b000001101010001111111101;
         rom[1975] = 24'b000001101001100001111011;
         rom[1976] = 24'b000001100100010110101110;
         rom[1977] = 24'b000001011111110100100010;
         rom[1978] = 24'b000001001011000011110101;
         rom[1979] = 24'b000001000101010111111000;
         rom[1980] = 24'b000001000001010100101111;
         rom[1981] = 24'b000000111010001111110111;
         rom[1982] = 24'b000000101111011111101111;
         rom[1983] = 24'b000000101001111010000110;
         rom[1984] = 24'b000000100110001101011000;
         rom[1985] = 24'b000000100010001011100111;
         rom[1986] = 24'b000000100001000111100101;
         rom[1987] = 24'b000000001111100110000010;
         rom[1988] = 24'b111111111011110101101101;
         rom[1989] = 24'b111111111101000101010100;
         rom[1990] = 24'b111111110100110001001101;
         rom[1991] = 24'b000000001100001010110001;
         rom[1992] = 24'b111111110110001111001010;
         rom[1993] = 24'b000000001101001000010100;
         rom[1994] = 24'b111111110110001110000111;
         rom[1995] = 24'b000000001000011001110011;
         rom[1996] = 24'b111111111100001001110111;
         rom[1997] = 24'b000000010000100111101100;
         rom[1998] = 24'b111111111111111111010100;
         rom[1999] = 24'b000000000001110101111110;
         end 

	 always @(posedge(clk))
		 begin 
			 if(reset) 
				 begin 
					 data_out <= 24'b0; 
					 i <= 16'b0; 
					 counter <= 16'b0; 
				 end 
			 else 
				 begin 
					 if(counter == 16'd5000) 
						 begin 
							 data_out <= rom[i]; 
							 counter <=16'b0; 
							 if(i == 1999) i <= 0; 
							 else i <= i + 1; 
						 end 
					 else counter <= counter + 16'd1; 
				 end 
		 end 

endmodule
