module gen_sinus( 
 	 output reg signed [23:0] data_out,
	 input clk,
	 input reset
	 ); 

	 reg signed [23:0] rom[0:39];
	 reg [15:0] i;
	 reg [15:0] counter;

	 always @(reset)
		 begin 
         rom[0] = 24'b000000000000000000000000;
         rom[1] = 24'b000011001000111001001001;
         rom[2] = 24'b000101011100011001101011;
         rom[3] = 24'b000110100010110101000101;
         rom[4] = 24'b000110101110100000011100;
         rom[5] = 24'b000110101111100101010111;
         rom[6] = 24'b000111010110011110001011;
         rom[7] = 24'b001000110110010001101010;
         rom[8] = 24'b001010111000100100110010;
         rom[9] = 24'b001100101001101110001010;
         rom[10] = 24'b001101010110011111100000;
         rom[11] = 24'b001100101001101110001010;
         rom[12] = 24'b001010111000100100110010;
         rom[13] = 24'b001000110110010001101010;
         rom[14] = 24'b000111010110011110001011;
         rom[15] = 24'b000110101111100101010111;
         rom[16] = 24'b000110101110100000011100;
         rom[17] = 24'b000110100010110101000101;
         rom[18] = 24'b000101011100011001101011;
         rom[19] = 24'b000011001000111001001001;
         rom[20] = 24'b000000000000000000000000;
         rom[21] = 24'b111100110111000110110111;
         rom[22] = 24'b111010100011100110010101;
         rom[23] = 24'b111001011101001010111011;
         rom[24] = 24'b111001010001011111100100;
         rom[25] = 24'b111001010000011010101001;
         rom[26] = 24'b111000101001100001110101;
         rom[27] = 24'b110111001001101110010110;
         rom[28] = 24'b110101000111011011001110;
         rom[29] = 24'b110011010110010001110110;
         rom[30] = 24'b110010101001100000100000;
         rom[31] = 24'b110011010110010001110110;
         rom[32] = 24'b110101000111011011001110;
         rom[33] = 24'b110111001001101110010110;
         rom[34] = 24'b111000101001100001110101;
         rom[35] = 24'b111001010000011010101001;
         rom[36] = 24'b111001010001011111100100;
         rom[37] = 24'b111001011101001010111011;
         rom[38] = 24'b111010100011100110010101;
         rom[39] = 24'b111100110111000110110111;
      end 

	 always @(posedge(clk))
		 begin 
			 if(reset) 
				 begin 
					 data_out <= 24'b0; 
					 i <= 16'b0; 
					 counter <= 16'b0; 
				 end 
			 else 
				 begin 
					 if(counter == 16'd5000) 
						 begin 
							 data_out <= rom[i]; 
							 counter <= 16'b0; 
							 if(i == 39) i <= 0; 
							 else i <= i + 1; 
						 end 
					 else counter <= counter + 16'd1; 
				 end 
		 end 

endmodule
