module gen_sinus( 
 	 output reg signed [23:0] data_out,
	 input clk,
	 input reset
	 ); 

	 reg signed [23:0] rom[0:39];
	 reg [15:0] i;
	 reg [15:0] counter;

	 always @(reset)
		 begin 
			 rom[0] = 24'b000000000000000000000000;
			 rom[1] = 24'b000001011111011110101110;
			 rom[2] = 24'b000010111100100110111110;
			 rom[3] = 24'b000100010101000110000000;
			 rom[4] = 24'b000101100110110000010111;
			 rom[5] = 24'b000110101111100101010111;
			 rom[6] = 24'b000111101101110010001110;
			 rom[7] = 24'b001000011111110100111100;
			 rom[8] = 24'b001001000100011110101001;
			 rom[9] = 24'b001001011010110101100101;
			 rom[10] = 24'b001001100010010110100000;
			 rom[11] = 24'b001001011010110101100101;
			 rom[12] = 24'b001001000100011110101001;
			 rom[13] = 24'b001000011111110100111100;
			 rom[14] = 24'b000111101101110010001110;
			 rom[15] = 24'b000110101111100101010111;
			 rom[16] = 24'b000101100110110000010111;
			 rom[17] = 24'b000100010101000110000000;
			 rom[18] = 24'b000010111100100110111110;
			 rom[19] = 24'b000001011111011110101110;
			 rom[20] = 24'b000000000000000000000000;
			 rom[21] = 24'b111110100000100001010010;
			 rom[22] = 24'b111101000011011001000010;
			 rom[23] = 24'b111011101010111010000000;
			 rom[24] = 24'b111010011001001111101001;
			 rom[25] = 24'b111001010000011010101001;
			 rom[26] = 24'b111000010010001101110010;
			 rom[27] = 24'b110111100000001011000100;
			 rom[28] = 24'b110110111011100001010111;
			 rom[29] = 24'b110110100101001010011011;
			 rom[30] = 24'b110110011101101001100000;
			 rom[31] = 24'b110110100101001010011011;
			 rom[32] = 24'b110110111011100001010111;
			 rom[33] = 24'b110111100000001011000100;
			 rom[34] = 24'b111000010010001101110010;
			 rom[35] = 24'b111001010000011010101001;
			 rom[36] = 24'b111010011001001111101001;
			 rom[37] = 24'b111011101010111010000000;
			 rom[38] = 24'b111101000011011001000010;
			 rom[39] = 24'b111110100000100001010010;
		 end 

	 always @(posedge(clk))
		 begin 
			 if(reset) 
				 begin 
					 data_out <= 24'b0; 
					 i <= 16'b0; 
					 counter <= 16'b0; 
				 end 
			 else 
				 begin 
					 if(counter == 16'd50000) 
						 begin 
							 data_out <= rom[i]; 
							 counter <= 16'b0; 
							 if(i == 39) i <= 0; 
							 else i <= i + 1; 
						 end 
					 else counter <= counter + 16'd1; 
				 end 
		 end 

endmodule
