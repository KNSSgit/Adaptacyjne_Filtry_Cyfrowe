module gen_ekg_50(
 	 output reg signed [23:0] data_out,
	 input clk,
	 input reset
	 ); 

	 reg signed [23:0] rom[0:1999];
	 reg [15:0] i;
	 reg [15:0] counter;//5000 * 2000pr�bek = 10 000 000 ; zegar 10mhz => 1hz

	 always @(reset)     // fs = 2kHz; f1 = 1Hz; A1 = 3000000; f2 = 50Hz; A2 = 90000
		 begin 
rom[0] = 24'b111111110101110110001110;
         rom[1] = 24'b000000000011001100001011;
         rom[2] = 24'b000000001101001100110000;
         rom[3] = 24'b000000001101011101001000;
         rom[4] = 24'b000000010110010101010010;
         rom[5] = 24'b000000001111000010011001;
         rom[6] = 24'b000000010010110000100001;
         rom[7] = 24'b000000100101101110100110;
         rom[8] = 24'b000000011101100100001000;
         rom[9] = 24'b000000011010101010000101;
         rom[10] = 24'b000000101100001011101111;
         rom[11] = 24'b000000101100000100110000;
         rom[12] = 24'b000000011111101111110110;
         rom[13] = 24'b000000100001011010001100;
         rom[14] = 24'b000000110000100011011010;
         rom[15] = 24'b000000010100010110010011;
         rom[16] = 24'b000000010100111101100001;
         rom[17] = 24'b000000010001011100010000;
         rom[18] = 24'b000000000111001101111110;
         rom[19] = 24'b000000001000011000000100;
         rom[20] = 24'b111111111000000101101101;
         rom[21] = 24'b111111110101101101010011;
         rom[22] = 24'b111111110110110111011011;
         rom[23] = 24'b111111011101110100111101;
         rom[24] = 24'b111111101110001111001011;
         rom[25] = 24'b111111100100100000001011;
         rom[26] = 24'b111111010110011111101001;
         rom[27] = 24'b111111011001101000101101;
         rom[28] = 24'b111111010011111111100000;
         rom[29] = 24'b111111011111101011101100;
         rom[30] = 24'b111111011111011110111100;
         rom[31] = 24'b111111100001100100001010;
         rom[32] = 24'b111111011101101111101001;
         rom[33] = 24'b111111100001011010110000;
         rom[34] = 24'b111111101011011001001010;
         rom[35] = 24'b111111011110101001011100;
         rom[36] = 24'b111111110010110000111011;
         rom[37] = 24'b111111101100011111000011;
         rom[38] = 24'b111111111001001101010110;
         rom[39] = 24'b111111110011101110011110;
         rom[40] = 24'b111111110110000011110111;
         rom[41] = 24'b000000001000111111110011;
         rom[42] = 24'b000000001000001101001100;
         rom[43] = 24'b000000001101011010011111;
         rom[44] = 24'b000000010110100100100011;
         rom[45] = 24'b000000100000111000010111;
         rom[46] = 24'b000000001111101010100101;
         rom[47] = 24'b000000011110110010101011;
         rom[48] = 24'b000000010010100010110100;
         rom[49] = 24'b000000110101001111010001;
         rom[50] = 24'b000000011111011111100000;
         rom[51] = 24'b000000100011111101100000;
         rom[52] = 24'b000000101101100001010110;
         rom[53] = 24'b000000011001000010110100;
         rom[54] = 24'b000000101000010101010010;
         rom[55] = 24'b000000011010111000000100;
         rom[56] = 24'b000000010110000111100001;
         rom[57] = 24'b000000010100011111000011;
         rom[58] = 24'b000000000101101010010100;
         rom[59] = 24'b000000010010000000010111;
         rom[60] = 24'b111111111010010100011100;
         rom[61] = 24'b111111110110100111001110;
         rom[62] = 24'b000000000000100000011110;
         rom[63] = 24'b111111100100000000011110;
         rom[64] = 24'b111111100111111010110010;
         rom[65] = 24'b111111101100010010101100;
         rom[66] = 24'b111111010010010110000001;
         rom[67] = 24'b111111011001011111001111;
         rom[68] = 24'b111111011101000011000010;
         rom[69] = 24'b111111011010101110111000;
         rom[70] = 24'b111111010100101001111100;
         rom[71] = 24'b111111101001101011001101;
         rom[72] = 24'b111111011011010100000101;
         rom[73] = 24'b111111100000011101111011;
         rom[74] = 24'b111111100101011101110110;
         rom[75] = 24'b111111101100100000110011;
         rom[76] = 24'b111111110001011011010111;
         rom[77] = 24'b111111110001001111101000;
         rom[78] = 24'b111111111101000011011111;
         rom[79] = 24'b111111111101110101011001;
         rom[80] = 24'b111111111100011001010111;
         rom[81] = 24'b000000000011001001010111;
         rom[82] = 24'b000000000101010010000111;
         rom[83] = 24'b000000011111110111100001;
         rom[84] = 24'b000000010101010110011010;
         rom[85] = 24'b000000011000001101010101;
         rom[86] = 24'b000000011010011111111100;
         rom[87] = 24'b000000100011001001110100;
         rom[88] = 24'b000000100101100001111111;
         rom[89] = 24'b000000110011110000010000;
         rom[90] = 24'b000000100000101101010110;
         rom[91] = 24'b000000100001010100110001;
         rom[92] = 24'b000000101000100110010111;
         rom[93] = 24'b000000011010010001001011;
         rom[94] = 24'b000000100000011001011110;
         rom[95] = 24'b000000010110001010101011;
         rom[96] = 24'b000000011010010011111110;
         rom[97] = 24'b000000100101100010000101;
         rom[98] = 24'b000000000111111000011110;
         rom[99] = 24'b000000000111011111110100;
         rom[100] = 24'b000000000110000010100110;
         rom[101] = 24'b111111111100101001001100;
         rom[102] = 24'b111111101001010011100010;
         rom[103] = 24'b111111100100010111110111;
         rom[104] = 24'b111111101100001100111010;
         rom[105] = 24'b111111011111011001110101;
         rom[106] = 24'b111111100000101110111010;
         rom[107] = 24'b111111011110011111001010;
         rom[108] = 24'b111111101101011011100111;
         rom[109] = 24'b111111110000100011111000;
         rom[110] = 24'b111111010110000000100100;
         rom[111] = 24'b111111001011000010011011;
         rom[112] = 24'b111111100111000110011111;
         rom[113] = 24'b111111001101110111101101;
         rom[114] = 24'b111111011010101100011110;
         rom[115] = 24'b111111101000000001100111;
         rom[116] = 24'b111111011101100001001110;
         rom[117] = 24'b111111111001011001010010;
         rom[118] = 24'b111111101010111110100110;
         rom[119] = 24'b111111111010111110111010;
         rom[120] = 24'b000000000010110001111101;
         rom[121] = 24'b111111110001110010010101;
         rom[122] = 24'b000000000001010010110111;
         rom[123] = 24'b000000000101110100110011;
         rom[124] = 24'b000000010011100010111111;
         rom[125] = 24'b000000010111011111111001;
         rom[126] = 24'b000000010101000000110010;
         rom[127] = 24'b000000011110100110100100;
         rom[128] = 24'b000000010100011010010101;
         rom[129] = 24'b000000100000001100010001;
         rom[130] = 24'b000000101000001010101000;
         rom[131] = 24'b000000101011000111101000;
         rom[132] = 24'b000000011111100110010100;
         rom[133] = 24'b000000101010101100100101;
         rom[134] = 24'b000000011001011100111000;
         rom[135] = 24'b000000011111000000000110;
         rom[136] = 24'b000000010101110100000001;
         rom[137] = 24'b000000001110001001111000;
         rom[138] = 24'b000000010000001011111011;
         rom[139] = 24'b000000000110100011100110;
         rom[140] = 24'b000000000110110011101010;
         rom[141] = 24'b000000000111010010110100;
         rom[142] = 24'b111111100101101101000011;
         rom[143] = 24'b111111111011111010111100;
         rom[144] = 24'b111111101010001010111101;
         rom[145] = 24'b111111100111000001111011;
         rom[146] = 24'b111111011100001110011010;
         rom[147] = 24'b111111011011010110100000;
         rom[148] = 24'b111111100001110011101001;
         rom[149] = 24'b111111010111001110000011;
         rom[150] = 24'b111111011001001110001001;
         rom[151] = 24'b111111011100100110110001;
         rom[152] = 24'b111111001011001101010111;
         rom[153] = 24'b111111100111100100001001;
         rom[154] = 24'b111111100110111011011001;
         rom[155] = 24'b111111011101011111110010;
         rom[156] = 24'b111111010101100111011001;
         rom[157] = 24'b111111110100011000010101;
         rom[158] = 24'b111111101100100111000101;
         rom[159] = 24'b111111110111100001001001;
         rom[160] = 24'b111111111100110001010000;
         rom[161] = 24'b111111110110010111100100;
         rom[162] = 24'b000000001010000000011011;
         rom[163] = 24'b000000001110010000000111;
         rom[164] = 24'b000000011010001100110001;
         rom[165] = 24'b000000010110110101100100;
         rom[166] = 24'b000000011010001110110011;
         rom[167] = 24'b000000011101110100111100;
         rom[168] = 24'b000000011100011111010000;
         rom[169] = 24'b000000100101111001101011;
         rom[170] = 24'b000000100011100010100000;
         rom[171] = 24'b000000011110100111100110;
         rom[172] = 24'b000000110011001100011100;
         rom[173] = 24'b000000100010001000111011;
         rom[174] = 24'b000000011010010000011101;
         rom[175] = 24'b000000011011110100001010;
         rom[176] = 24'b000000100000011011011100;
         rom[177] = 24'b000000000110111011110011;
         rom[178] = 24'b111111111100001101100100;
         rom[179] = 24'b000000001010111100001111;
         rom[180] = 24'b111111111010101110100000;
         rom[181] = 24'b000000000001110111001000;
         rom[182] = 24'b111111100111110110000101;
         rom[183] = 24'b111111101010010010011100;
         rom[184] = 24'b111111101111110011110010;
         rom[185] = 24'b111111100000100001010011;
         rom[186] = 24'b111111011101011011100100;
         rom[187] = 24'b111111011011111011011000;
         rom[188] = 24'b111111100100100001010110;
         rom[189] = 24'b111111010111010101110011;
         rom[190] = 24'b111111010101011000110110;
         rom[191] = 24'b111111011001000001101010;
         rom[192] = 24'b111111011101001100001101;
         rom[193] = 24'b111111011101010111101011;
         rom[194] = 24'b111111101000000111011100;
         rom[195] = 24'b111111100011001010110111;
         rom[196] = 24'b111111101010101001001111;
         rom[197] = 24'b111111101011111001010110;
         rom[198] = 24'b111111111100000100100111;
         rom[199] = 24'b000000000001101110001010;
         rom[200] = 24'b000000001001100101101011;
         rom[201] = 24'b000000000001100101001110;
         rom[202] = 24'b000000001000010100010110;
         rom[203] = 24'b000000100000010101100100;
         rom[204] = 24'b000000001111011011000101;
         rom[205] = 24'b000000001110110111011011;
         rom[206] = 24'b000000011001111101101101;
         rom[207] = 24'b000000100110101100010110;
         rom[208] = 24'b000000010111000001100110;
         rom[209] = 24'b000000100100111110101001;
         rom[210] = 24'b000000011111111010011101;
         rom[211] = 24'b000000101101001100100110;
         rom[212] = 24'b000000011101011110100000;
         rom[213] = 24'b000000010100100100001010;
         rom[214] = 24'b000000100100011100111011;
         rom[215] = 24'b000000101000101111011001;
         rom[216] = 24'b000000010001101101001111;
         rom[217] = 24'b000000001010001001001110;
         rom[218] = 24'b000000010110000000011110;
         rom[219] = 24'b111111111010011011101100;
         rom[220] = 24'b000000001000110011110001;
         rom[221] = 24'b111111110001011100100110;
         rom[222] = 24'b000000000111111100011000;
         rom[223] = 24'b111111100011011000010101;
         rom[224] = 24'b111111101011110111111111;
         rom[225] = 24'b111111100100010100011101;
         rom[226] = 24'b111111011110101001001101;
         rom[227] = 24'b111111011101010011110000;
         rom[228] = 24'b111111100100011010101011;
         rom[229] = 24'b111111010111110010111010;
         rom[230] = 24'b111111100001001010110011;
         rom[231] = 24'b111111100110000011110110;
         rom[232] = 24'b111111011101110111101101;
         rom[233] = 24'b111111100000110110011101;
         rom[234] = 24'b111111011101000100001011;
         rom[235] = 24'b111111101000101101000001;
         rom[236] = 24'b111111100010001110100110;
         rom[237] = 24'b111111110111100100111010;
         rom[238] = 24'b111111101100110101011011;
         rom[239] = 24'b111111110100000001010101;
         rom[240] = 24'b000000000101100011010100;
         rom[241] = 24'b000000000101010011010010;
         rom[242] = 24'b000000001001110100011010;
         rom[243] = 24'b000000010010110100111111;
         rom[244] = 24'b000000010110011001110101;
         rom[245] = 24'b000000010000101010110001;
         rom[246] = 24'b000000101001110101111011;
         rom[247] = 24'b000000010101001101010111;
         rom[248] = 24'b000000100111101000011010;
         rom[249] = 24'b000000101001000000100011;
         rom[250] = 24'b000000100011110010100000;
         rom[251] = 24'b000000100001101100011000;
         rom[252] = 24'b000000011101111010110100;
         rom[253] = 24'b000000001011000110111011;
         rom[254] = 24'b000000101001011111100011;
         rom[255] = 24'b000000011101100101101010;
         rom[256] = 24'b000000011100000011100100;
         rom[257] = 24'b000000001001110001010100;
         rom[258] = 24'b000000011010101101010001;
         rom[259] = 24'b000000001111100110101110;
         rom[260] = 24'b000000001001101100100001;
         rom[261] = 24'b111111111010000010001100;
         rom[262] = 24'b111111110011011110101100;
         rom[263] = 24'b111111110101011000011001;
         rom[264] = 24'b111111100111011011100101;
         rom[265] = 24'b111111100101100000010101;
         rom[266] = 24'b111111011100100000000111;
         rom[267] = 24'b111111011000011100111000;
         rom[268] = 24'b111111010111011000000000;
         rom[269] = 24'b111111011101110001101100;
         rom[270] = 24'b111111100010110010010110;
         rom[271] = 24'b111111100000001110111001;
         rom[272] = 24'b111111100001000011000010;
         rom[273] = 24'b111111010101110110001000;
         rom[274] = 24'b111111100111011001111010;
         rom[275] = 24'b111111101000000011000001;
         rom[276] = 24'b111111110101111101111001;
         rom[277] = 24'b111111101011111010000100;
         rom[278] = 24'b000000000110010011001011;
         rom[279] = 24'b000000001000111110001010;
         rom[280] = 24'b000000000010010010010110;
         rom[281] = 24'b000000000010101101101101;
         rom[282] = 24'b000000010011100111101111;
         rom[283] = 24'b000000010011011111110010;
         rom[284] = 24'b000000001011011000011010;
         rom[285] = 24'b000000011010000100100001;
         rom[286] = 24'b000000100111110110111111;
         rom[287] = 24'b000000011011101111010000;
         rom[288] = 24'b000000101101001000100010;
         rom[289] = 24'b000000101000011010010111;
         rom[290] = 24'b000000110100001110001101;
         rom[291] = 24'b000000100000001001101010;
         rom[292] = 24'b000000101001110001001101;
         rom[293] = 24'b000000100001100011110010;
         rom[294] = 24'b000000001100011110101111;
         rom[295] = 24'b000000011011001101001101;
         rom[296] = 24'b000000011000111111000010;
         rom[297] = 24'b000000010100110000101111;
         rom[298] = 24'b000000001101110111100011;
         rom[299] = 24'b000000000101101000111101;
         rom[300] = 24'b000000000000000011100111;
         rom[301] = 24'b111111111100001101100101;
         rom[302] = 24'b111111110010100000010101;
         rom[303] = 24'b111111110100100001010110;
         rom[304] = 24'b111111100111100111010100;
         rom[305] = 24'b111111100110110000111001;
         rom[306] = 24'b111111101000000101010001;
         rom[307] = 24'b111111011000110010010011;
         rom[308] = 24'b111111011110000011111111;
         rom[309] = 24'b111111001000101001101010;
         rom[310] = 24'b111111011000001000001010;
         rom[311] = 24'b111111010111000110111000;
         rom[312] = 24'b111111011100110100001100;
         rom[313] = 24'b111111011010011010110110;
         rom[314] = 24'b111111011111111011111111;
         rom[315] = 24'b111111100010010101101001;
         rom[316] = 24'b111111101001100111000011;
         rom[317] = 24'b111111111110100110111010;
         rom[318] = 24'b111111110001100111011110;
         rom[319] = 24'b000000000001101000000011;
         rom[320] = 24'b111111110111110101010000;
         rom[321] = 24'b000000001110110110100010;
         rom[322] = 24'b000000000010001101001110;
         rom[323] = 24'b000000010111000110101010;
         rom[324] = 24'b000000001111001100100001;
         rom[325] = 24'b000000010111011100000101;
         rom[326] = 24'b000000011101000001011000;
         rom[327] = 24'b000000100001001010100010;
         rom[328] = 24'b000000010111001110111101;
         rom[329] = 24'b000000101000000010000001;
         rom[330] = 24'b000000101100101001100011;
         rom[331] = 24'b000000011111001101011001;
         rom[332] = 24'b000000011101111100111000;
         rom[333] = 24'b000000100101110100000101;
         rom[334] = 24'b000000100000100011110010;
         rom[335] = 24'b000000010111101111011101;
         rom[336] = 24'b000000010100010001010100;
         rom[337] = 24'b000000011110010111100110;
         rom[338] = 24'b000000000101010010111100;
         rom[339] = 24'b000000000110110101111000;
         rom[340] = 24'b000000000001000000010100;
         rom[341] = 24'b111111111110101111010110;
         rom[342] = 24'b111111111111101010110101;
         rom[343] = 24'b111111101010110100000010;
         rom[344] = 24'b111111100101101110010101;
         rom[345] = 24'b111111011100100011111100;
         rom[346] = 24'b111111010111111010101011;
         rom[347] = 24'b111111010110100110000111;
         rom[348] = 24'b111111011000110001111011;
         rom[349] = 24'b111111011010100011000010;
         rom[350] = 24'b111111100010101011110101;
         rom[351] = 24'b111111010000100101101001;
         rom[352] = 24'b111111100010100110101001;
         rom[353] = 24'b111111100101111001010011;
         rom[354] = 24'b111111100001101010101101;
         rom[355] = 24'b111111100001110010001011;
         rom[356] = 24'b111111110010001000100110;
         rom[357] = 24'b111111101001100111101001;
         rom[358] = 24'b111111111001100101100011;
         rom[359] = 24'b111111111000010101101010;
         rom[360] = 24'b111111111101110011101110;
         rom[361] = 24'b000000000010000110100000;
         rom[362] = 24'b000000000001001011110100;
         rom[363] = 24'b000000010001111000010000;
         rom[364] = 24'b000000011100101001010110;
         rom[365] = 24'b000000011111111101111101;
         rom[366] = 24'b000000011100110111011110;
         rom[367] = 24'b000000101001001111011110;
         rom[368] = 24'b000000010000111111001010;
         rom[369] = 24'b000000100001010100111110;
         rom[370] = 24'b000000100001101011011111;
         rom[371] = 24'b000000110100001101110111;
         rom[372] = 24'b000000100100011110100001;
         rom[373] = 24'b000000010110101110111011;
         rom[374] = 24'b000000100001100001100100;
         rom[375] = 24'b000000011101111010101000;
         rom[376] = 24'b000000001111011001001010;
         rom[377] = 24'b000000011001000110011110;
         rom[378] = 24'b000000001100011011000110;
         rom[379] = 24'b000000001011101000100010;
         rom[380] = 24'b111111111111111100101010;
         rom[381] = 24'b000000000101101110110011;
         rom[382] = 24'b111111111000001110010110;
         rom[383] = 24'b111111101110100100010111;
         rom[384] = 24'b111111100111110001000001;
         rom[385] = 24'b111111101000110111110010;
         rom[386] = 24'b111111100110000010100111;
         rom[387] = 24'b111111010101001111010001;
         rom[388] = 24'b111111100001101100001000;
         rom[389] = 24'b111111011100001100000110;
         rom[390] = 24'b111111100001100000010000;
         rom[391] = 24'b111111011011111110000001;
         rom[392] = 24'b111111100100000001010011;
         rom[393] = 24'b111111100100111100011010;
         rom[394] = 24'b111111101011001010110011;
         rom[395] = 24'b111111100011011111011010;
         rom[396] = 24'b111111111001010100000101;
         rom[397] = 24'b111111100111010010010010;
         rom[398] = 24'b111111111111100011011000;
         rom[399] = 24'b000000000011100000110100;
         rom[400] = 24'b000000000001000101110011;
         rom[401] = 24'b000000000000100011010101;
         rom[402] = 24'b000000010001110110100111;
         rom[403] = 24'b111111111111101010010000;
         rom[404] = 24'b000000011111101011111101;
         rom[405] = 24'b000000011110000000000000;
         rom[406] = 24'b000000010011010111101111;
         rom[407] = 24'b000000100100011011101101;
         rom[408] = 24'b000000101100000000001111;
         rom[409] = 24'b000000010010110011001111;
         rom[410] = 24'b000000100111100000110010;
         rom[411] = 24'b000000011111111111000000;
         rom[412] = 24'b000000100101001000010010;
         rom[413] = 24'b000000100100010010101100;
         rom[414] = 24'b000000011000111001001111;
         rom[415] = 24'b000000010111010100110110;
         rom[416] = 24'b000000010010101001101001;
         rom[417] = 24'b000000001000011000001100;
         rom[418] = 24'b000000010100011111000110;
         rom[419] = 24'b111111110010110101011110;
         rom[420] = 24'b111111111000000000110010;
         rom[421] = 24'b111111110110111110111101;
         rom[422] = 24'b111111111101101011010010;
         rom[423] = 24'b111111101110010110101110;
         rom[424] = 24'b111111101011000000101111;
         rom[425] = 24'b111111100111010010001100;
         rom[426] = 24'b111111011100001001001001;
         rom[427] = 24'b111111100001010000111010;
         rom[428] = 24'b111111100011100011100001;
         rom[429] = 24'b111111011101101011011100;
         rom[430] = 24'b111111001100001010010110;
         rom[431] = 24'b111111011010000101001110;
         rom[432] = 24'b111111011001101111100100;
         rom[433] = 24'b111111100100111100001110;
         rom[434] = 24'b111111011101000110000000;
         rom[435] = 24'b111111100111110111111100;
         rom[436] = 24'b111111100110100110011111;
         rom[437] = 24'b111111100100011001110010;
         rom[438] = 24'b111111110101110010001111;
         rom[439] = 24'b000000000001000100000011;
         rom[440] = 24'b000000000011111011001000;
         rom[441] = 24'b000000000011011111101001;
         rom[442] = 24'b000000000110110101010111;
         rom[443] = 24'b111111111111101110001011;
         rom[444] = 24'b000000011001000010110011;
         rom[445] = 24'b000000010101111011111111;
         rom[446] = 24'b000000010010101010110000;
         rom[447] = 24'b000000100000111111110110;
         rom[448] = 24'b000000100011110001100001;
         rom[449] = 24'b000000110001111100100011;
         rom[450] = 24'b000000011001000111101001;
         rom[451] = 24'b000000101001000000000111;
         rom[452] = 24'b000000100100101000001011;
         rom[453] = 24'b000000100101001101000110;
         rom[454] = 24'b000000100011011000100100;
         rom[455] = 24'b000000100101001001110111;
         rom[456] = 24'b000000000111000011100110;
         rom[457] = 24'b000000000110111011010100;
         rom[458] = 24'b000000000111000111100100;
         rom[459] = 24'b111111111010101101100001;
         rom[460] = 24'b111111110001100100111000;
         rom[461] = 24'b111111111100111101100110;
         rom[462] = 24'b111111111111010101000110;
         rom[463] = 24'b111111110001110010010011;
         rom[464] = 24'b111111011010000110101111;
         rom[465] = 24'b111111011111001110001000;
         rom[466] = 24'b111111100010001000010111;
         rom[467] = 24'b111111010011010001001001;
         rom[468] = 24'b111111101000011011000001;
         rom[469] = 24'b111111011110110101010100;
         rom[470] = 24'b111111011100111111111001;
         rom[471] = 24'b111111011001111100110110;
         rom[472] = 24'b111111100011000011111011;
         rom[473] = 24'b111111100010010001001111;
         rom[474] = 24'b111111011101101101100011;
         rom[475] = 24'b111111100100000011000101;
         rom[476] = 24'b111111111010101001011001;
         rom[477] = 24'b111111101000000000011010;
         rom[478] = 24'b111111111001101110100011;
         rom[479] = 24'b000000001000011011101110;
         rom[480] = 24'b111111111100111101111110;
         rom[481] = 24'b000000001011010000100111;
         rom[482] = 24'b000000011110101000101010;
         rom[483] = 24'b000000000111101010110100;
         rom[484] = 24'b000000001111111100100111;
         rom[485] = 24'b000000100101101101001101;
         rom[486] = 24'b000000101000100011110001;
         rom[487] = 24'b000000011110111011000110;
         rom[488] = 24'b000000100000101100111100;
         rom[489] = 24'b000000011000000101001000;
         rom[490] = 24'b000000101010110101111001;
         rom[491] = 24'b000000110001001101011111;
         rom[492] = 24'b000000100100110100001110;
         rom[493] = 24'b000000011010010101010001;
         rom[494] = 24'b000000011100011111111000;
         rom[495] = 24'b000000010100010010001000;
         rom[496] = 24'b000000010101010111101110;
         rom[497] = 24'b000000010001001000000000;
         rom[498] = 24'b000000001111101111001001;
         rom[499] = 24'b111111111000100111100010;
         rom[500] = 24'b000000001010000111000011;
         rom[501] = 24'b111111111001010100000100;
         rom[502] = 24'b111111101111101010100111;
         rom[503] = 24'b111111110000111111000111;
         rom[504] = 24'b111111100100101001011111;
         rom[505] = 24'b111111100001110001010110;
         rom[506] = 24'b111111011110111101001000;
         rom[507] = 24'b111111010011111101111001;
         rom[508] = 24'b111111011001100010000001;
         rom[509] = 24'b111111100011011001110011;
         rom[510] = 24'b111111100111010101010001;
         rom[511] = 24'b111111011011110100100101;
         rom[512] = 24'b111111100010001100100110;
         rom[513] = 24'b111111011111001011001000;
         rom[514] = 24'b111111010110000000100101;
         rom[515] = 24'b111111100101010110110110;
         rom[516] = 24'b111111110101000110010100;
         rom[517] = 24'b111111110001100001010110;
         rom[518] = 24'b111111111000000110010100;
         rom[519] = 24'b111111110011110110010111;
         rom[520] = 24'b111111110011111100100000;
         rom[521] = 24'b000000000101100001010110;
         rom[522] = 24'b000000001001100100110000;
         rom[523] = 24'b000000000101001000000101;
         rom[524] = 24'b000000001001000100100111;
         rom[525] = 24'b000000010101011001000101;
         rom[526] = 24'b000000100000011001111111;
         rom[527] = 24'b000000100011000100001100;
         rom[528] = 24'b000000101010101010111100;
         rom[529] = 24'b000000011100010110001111;
         rom[530] = 24'b000000100011101000001111;
         rom[531] = 24'b000000011000111111100100;
         rom[532] = 24'b000000100000110000100100;
         rom[533] = 24'b000000010011100011011000;
         rom[534] = 24'b000000101000100001010010;
         rom[535] = 24'b000000010110110110001110;
         rom[536] = 24'b000000010011010111110110;
         rom[537] = 24'b000000010110100110100010;
         rom[538] = 24'b000000000110011101000000;
         rom[539] = 24'b000000000100001110001000;
         rom[540] = 24'b111111111101110100010000;
         rom[541] = 24'b111111111011001110001101;
         rom[542] = 24'b111111110011010001111110;
         rom[543] = 24'b111111111111010010101110;
         rom[544] = 24'b111111101001000010011101;
         rom[545] = 24'b111111100111111000001101;
         rom[546] = 24'b111111100111000111110000;
         rom[547] = 24'b111111011101100110100001;
         rom[548] = 24'b111111100111101100110001;
         rom[549] = 24'b111111010111111000000101;
         rom[550] = 24'b111111001010001001101100;
         rom[551] = 24'b111111011100101101101111;
         rom[552] = 24'b111111011010011010000011;
         rom[553] = 24'b111111011110100111010001;
         rom[554] = 24'b111111110000101010110010;
         rom[555] = 24'b111111101100000100111111;
         rom[556] = 24'b111111101011000101111111;
         rom[557] = 24'b111111111010010101110111;
         rom[558] = 24'b111111110001101010010100;
         rom[559] = 24'b111111111100001010100100;
         rom[560] = 24'b111111111111010100011111;
         rom[561] = 24'b000000010110111100100011;
         rom[562] = 24'b000000001111110100100101;
         rom[563] = 24'b000000010001110100011000;
         rom[564] = 24'b000000001010111100100110;
         rom[565] = 24'b000000010111110001001100;
         rom[566] = 24'b000000010100100001010000;
         rom[567] = 24'b000000100111110001001110;
         rom[568] = 24'b000000011111111011111010;
         rom[569] = 24'b000000010110101011001110;
         rom[570] = 24'b000000011100111011111010;
         rom[571] = 24'b000000100111101000111010;
         rom[572] = 24'b000000011101111000000010;
         rom[573] = 24'b000000100011000111110011;
         rom[574] = 24'b000000101011100111110110;
         rom[575] = 24'b000000100000101101010111;
         rom[576] = 24'b000000100011110011000010;
         rom[577] = 24'b000000001100011101010000;
         rom[578] = 24'b000000001110001110110101;
         rom[579] = 24'b111111111110111100111010;
         rom[580] = 24'b111111111110111100101010;
         rom[581] = 24'b111111111011011000000111;
         rom[582] = 24'b111111110010011010101011;
         rom[583] = 24'b111111111000111101111011;
         rom[584] = 24'b111111110110010000010100;
         rom[585] = 24'b111111101000100101100111;
         rom[586] = 24'b111111011111011011101100;
         rom[587] = 24'b111111011110010111100110;
         rom[588] = 24'b111111010110001100000111;
         rom[589] = 24'b111111011001100000100101;
         rom[590] = 24'b111111011000110101000100;
         rom[591] = 24'b111111100101100100000001;
         rom[592] = 24'b111111011001101100110100;
         rom[593] = 24'b111111011100111000000010;
         rom[594] = 24'b111111101101110001000111;
         rom[595] = 24'b111111011011010101101111;
         rom[596] = 24'b111111100111110011101101;
         rom[597] = 24'b111111110001011011001011;
         rom[598] = 24'b111111110000001000010000;
         rom[599] = 24'b000000000011001001011010;
         rom[600] = 24'b111111111001110110110110;
         rom[601] = 24'b000000000011010011111000;
         rom[602] = 24'b111111111101011000001100;
         rom[603] = 24'b000000001111011001000000;
         rom[604] = 24'b000000011111111111100001;
         rom[605] = 24'b000000010111111010111010;
         rom[606] = 24'b000000101011100000011101;
         rom[607] = 24'b000000011111011111001001;
         rom[608] = 24'b000000010100111101001011;
         rom[609] = 24'b000000100101001100101001;
         rom[610] = 24'b000000101001110000000011;
         rom[611] = 24'b000000100100011110110001;
         rom[612] = 24'b000000100010100001100011;
         rom[613] = 24'b000000011111100000010010;
         rom[614] = 24'b000000101001011010110001;
         rom[615] = 24'b000000011010101101001011;
         rom[616] = 24'b000000010101000111110010;
         rom[617] = 24'b000000011110100100111000;
         rom[618] = 24'b000000000011111111000000;
         rom[619] = 24'b111111111001110100101000;
         rom[620] = 24'b000000000101111000110001;
         rom[621] = 24'b111111111010100011000101;
         rom[622] = 24'b111111110110111111011011;
         rom[623] = 24'b111111110000101100000100;
         rom[624] = 24'b111111101001101111110101;
         rom[625] = 24'b111111100101100000101100;
         rom[626] = 24'b111111010010011010011101;
         rom[627] = 24'b111111010100001101010001;
         rom[628] = 24'b111111100000111010000100;
         rom[629] = 24'b111111100110100010001111;
         rom[630] = 24'b111111010010001010011110;
         rom[631] = 24'b111111010000101101101011;
         rom[632] = 24'b111111100101000101100100;
         rom[633] = 24'b111111011111010111010010;
         rom[634] = 24'b111111011111100110010101;
         rom[635] = 24'b111111100110101101111110;
         rom[636] = 24'b111111110001010111101001;
         rom[637] = 24'b111111101101110111110100;
         rom[638] = 24'b111111101100011001011000;
         rom[639] = 24'b000000000110100100101100;
         rom[640] = 24'b111111111011100100001011;
         rom[641] = 24'b111111111100011000011011;
         rom[642] = 24'b000000001000010111100110;
         rom[643] = 24'b000000010101110111001000;
         rom[644] = 24'b000000001110001100010011;
         rom[645] = 24'b000000011001110111010110;
         rom[646] = 24'b000000011110000010101111;
         rom[647] = 24'b000000100011001101101111;
         rom[648] = 24'b000000011100001111101101;
         rom[649] = 24'b000000100000101001100101;
         rom[650] = 24'b000000011110011110010000;
         rom[651] = 24'b000000100100101010101110;
         rom[652] = 24'b000000101111100111111101;
         rom[653] = 24'b000000101000010001110010;
         rom[654] = 24'b000000101111010101010110;
         rom[655] = 24'b000000011010010110011100;
         rom[656] = 24'b000000010110011001101001;
         rom[657] = 24'b000000001101101000011110;
         rom[658] = 24'b000000001000100110011000;
         rom[659] = 24'b000000000110000101010110;
         rom[660] = 24'b000000000000111000000111;
         rom[661] = 24'b111111110101011110101110;
         rom[662] = 24'b111111110110101000110000;
         rom[663] = 24'b111111110010011000101111;
         rom[664] = 24'b111111101101000100101110;
         rom[665] = 24'b111111100101100010001110;
         rom[666] = 24'b111111101010001010100111;
         rom[667] = 24'b111111011111000111111011;
         rom[668] = 24'b111111011100011111001010;
         rom[669] = 24'b111111001111111010001111;
         rom[670] = 24'b111111011001000010100011;
         rom[671] = 24'b111111101011010000011010;
         rom[672] = 24'b111111100101010011100110;
         rom[673] = 24'b111111001110111110000011;
         rom[674] = 24'b111111101011101011010011;
         rom[675] = 24'b111111101011000111100000;
         rom[676] = 24'b111111100010011110000111;
         rom[677] = 24'b111111110000110010001110;
         rom[678] = 24'b111111110110101110000000;
         rom[679] = 24'b000000000110011010100100;
         rom[680] = 24'b111111111011100101101101;
         rom[681] = 24'b111111111101110000000101;
         rom[682] = 24'b000000001111110100010000;
         rom[683] = 24'b000000010111000001110101;
         rom[684] = 24'b000000010001111000010111;
         rom[685] = 24'b000000100011100000010000;
         rom[686] = 24'b000000011011000001111010;
         rom[687] = 24'b000000011111001010100100;
         rom[688] = 24'b000000011001000111011100;
         rom[689] = 24'b000000101011110011010110;
         rom[690] = 24'b000000101011011110001111;
         rom[691] = 24'b000000100101011010000001;
         rom[692] = 24'b000000010100101011101101;
         rom[693] = 24'b000000101000111110110001;
         rom[694] = 24'b000000100011001000100101;
         rom[695] = 24'b000000011000001010110001;
         rom[696] = 24'b000000010000100010001110;
         rom[697] = 24'b000000001010100010010101;
         rom[698] = 24'b000000000000000110111000;
         rom[699] = 24'b111111111000001011101000;
         rom[700] = 24'b111111111111100110101011;
         rom[701] = 24'b111111110100000101100001;
         rom[702] = 24'b111111110111100000110110;
         rom[703] = 24'b111111110010101110101001;
         rom[704] = 24'b111111100111110011010010;
         rom[705] = 24'b111111100111011011000111;
         rom[706] = 24'b111111101000001101001001;
         rom[707] = 24'b111111100000100110011110;
         rom[708] = 24'b111111100110000111110110;
         rom[709] = 24'b111111011100000101101010;
         rom[710] = 24'b111111010111000111110101;
         rom[711] = 24'b111111010011101010010001;
         rom[712] = 24'b111111010010000011110000;
         rom[713] = 24'b111111100100011111010100;
         rom[714] = 24'b111111101011101101101010;
         rom[715] = 24'b111111110001101000100101;
         rom[716] = 24'b111111100101011101011110;
         rom[717] = 24'b111111110100100110101001;
         rom[718] = 24'b111111101101100010010010;
         rom[719] = 24'b000000000000110110110101;
         rom[720] = 24'b111111111101010110010011;
         rom[721] = 24'b000000010101000001010000;
         rom[722] = 24'b000000010000101010111001;
         rom[723] = 24'b000000001100010010000000;
         rom[724] = 24'b000000100010000101011011;
         rom[725] = 24'b000000011110101011111100;
         rom[726] = 24'b000000100111101000110111;
         rom[727] = 24'b000000011100111111001110;
         rom[728] = 24'b000000101011011101011111;
         rom[729] = 24'b000000110000110110101011;
         rom[730] = 24'b000000100000101011011110;
         rom[731] = 24'b000000011110011001001111;
         rom[732] = 24'b000000101011101000010001;
         rom[733] = 24'b000000011100001110101000;
         rom[734] = 24'b000000100000010010011101;
         rom[735] = 24'b000000010101100101000001;
         rom[736] = 24'b000000010111001110110100;
         rom[737] = 24'b000000010100100111101100;
         rom[738] = 24'b000000010000000000001100;
         rom[739] = 24'b111111110111101001010100;
         rom[740] = 24'b111111110101101101101010;
         rom[741] = 24'b111111110000100011110110;
         rom[742] = 24'b111111111001110011000101;
         rom[743] = 24'b111111110101000001011001;
         rom[744] = 24'b111111100110110100001001;
         rom[745] = 24'b111111101010100101110001;
         rom[746] = 24'b111111101100100110000001;
         rom[747] = 24'b111111011101110111011001;
         rom[748] = 24'b111111011100101111100000;
         rom[749] = 24'b111111011010110000000110;
         rom[750] = 24'b111111010001101011001111;
         rom[751] = 24'b111111011111011001010010;
         rom[752] = 24'b111111001101000110011011;
         rom[753] = 24'b111111101010010101010011;
         rom[754] = 24'b111111101110001011101011;
         rom[755] = 24'b111111101011100100101110;
         rom[756] = 24'b111111110000001010111111;
         rom[757] = 24'b111111110001101010000100;
         rom[758] = 24'b000000000110101110001111;
         rom[759] = 24'b111111111000010101001001;
         rom[760] = 24'b111111110111000101100101;
         rom[761] = 24'b000000010001101110011101;
         rom[762] = 24'b000000000110010010010101;
         rom[763] = 24'b000000010111010100000011;
         rom[764] = 24'b000000001010110101110110;
         rom[765] = 24'b000000010001001010000011;
         rom[766] = 24'b000000100101000000001100;
         rom[767] = 24'b000000011111100000110010;
         rom[768] = 24'b000000101001011000000010;
         rom[769] = 24'b000000100100111111010110;
         rom[770] = 24'b000000101101010000101110;
         rom[771] = 24'b000000110010110101101111;
         rom[772] = 24'b000000011010110101011110;
         rom[773] = 24'b000000100110101001111100;
         rom[774] = 24'b000000011001100101011010;
         rom[775] = 24'b000000011100101110011001;
         rom[776] = 24'b000000010011010001100101;
         rom[777] = 24'b000000010100000100111101;
         rom[778] = 24'b000000001110001010011000;
         rom[779] = 24'b000000001000010010100010;
         rom[780] = 24'b111111110110001001001100;
         rom[781] = 24'b111111101110111111111100;
         rom[782] = 24'b111111111100111111100010;
         rom[783] = 24'b111111110001100100111011;
         rom[784] = 24'b111111100111011010000001;
         rom[785] = 24'b111111110101000111101010;
         rom[786] = 24'b111111100111001101010100;
         rom[787] = 24'b111111101100000000101111;
         rom[788] = 24'b111111011111000011111100;
         rom[789] = 24'b111111011011011011101101;
         rom[790] = 24'b111111011011101101000100;
         rom[791] = 24'b111111010011001000100100;
         rom[792] = 24'b111111100010101001000011;
         rom[793] = 24'b111111011111101101011100;
         rom[794] = 24'b111111100011000010101011;
         rom[795] = 24'b111111110101000111010001;
         rom[796] = 24'b111111110101110010111010;
         rom[797] = 24'b111111110011011101100111;
         rom[798] = 24'b111111110110001011010000;
         rom[799] = 24'b000000000111001111000101;
         rom[800] = 24'b111111111011011000101001;
         rom[801] = 24'b000000001000001010111100;
         rom[802] = 24'b000000000010110010111110;
         rom[803] = 24'b000000011011001100111011;
         rom[804] = 24'b000000011111011001110100;
         rom[805] = 24'b000000010101111101001011;
         rom[806] = 24'b000000010111001111110010;
         rom[807] = 24'b000000100101000110011010;
         rom[808] = 24'b000000101010010100001111;
         rom[809] = 24'b000000100000011111010101;
         rom[810] = 24'b000000010111111100100011;
         rom[811] = 24'b000000100101011011101000;
         rom[812] = 24'b000000011111010100011010;
         rom[813] = 24'b000000011011011000100110;
         rom[814] = 24'b000000010111101111100101;
         rom[815] = 24'b000000011101111001001110;
         rom[816] = 24'b000000011011000000111001;
         rom[817] = 24'b000000001100001100110001;
         rom[818] = 24'b000000000001001011011111;
         rom[819] = 24'b000000000000000111111001;
         rom[820] = 24'b000000000011101110000011;
         rom[821] = 24'b111111110101011100111110;
         rom[822] = 24'b111111111101110000000100;
         rom[823] = 24'b111111101111000000110111;
         rom[824] = 24'b111111101111100010011110;
         rom[825] = 24'b111111100101111110111110;
         rom[826] = 24'b111111100110000111001111;
         rom[827] = 24'b111111010011000100000101;
         rom[828] = 24'b111111100101010001010101;
         rom[829] = 24'b111111011100011101101000;
         rom[830] = 24'b111111100000100110011010;
         rom[831] = 24'b111111010011101010000100;
         rom[832] = 24'b111111100010111111101111;
         rom[833] = 24'b111111100101110110100000;
         rom[834] = 24'b111111011011010011000011;
         rom[835] = 24'b111111100100100010101111;
         rom[836] = 24'b111111101010001111010111;
         rom[837] = 24'b111111101100100111000101;
         rom[838] = 24'b111111111111100100011100;
         rom[839] = 24'b111111111011100110110100;
         rom[840] = 24'b000000000101100100100100;
         rom[841] = 24'b000000000010101000000111;
         rom[842] = 24'b000000010111111000011010;
         rom[843] = 24'b000000010011011010000101;
         rom[844] = 24'b000000010101111110000001;
         rom[845] = 24'b000000011010011110001001;
         rom[846] = 24'b000000011111101010111011;
         rom[847] = 24'b000000010110100001000100;
         rom[848] = 24'b000000101000000011001011;
         rom[849] = 24'b000000011100100101111100;
         rom[850] = 24'b000000100101001000111000;
         rom[851] = 24'b000000101001011101100010;
         rom[852] = 24'b000000011110010100100111;
         rom[853] = 24'b000000011111001101100011;
         rom[854] = 24'b000000010101101100111011;
         rom[855] = 24'b000000011011010101010100;
         rom[856] = 24'b000000011101101010101001;
         rom[857] = 24'b000000010110000100000001;
         rom[858] = 24'b000000000111000111011010;
         rom[859] = 24'b000000000101101101011100;
         rom[860] = 24'b111111111101100100000010;
         rom[861] = 24'b111111110100011101001011;
         rom[862] = 24'b111111110111010111011000;
         rom[863] = 24'b111111111000101010111101;
         rom[864] = 24'b111111101001101101010100;
         rom[865] = 24'b111111011111010011101111;
         rom[866] = 24'b111111100101010101100001;
         rom[867] = 24'b111111100010100010110001;
         rom[868] = 24'b111111100010011000010100;
         rom[869] = 24'b111111010101110001010010;
         rom[870] = 24'b111111011011111110101011;
         rom[871] = 24'b111111010011111010011000;
         rom[872] = 24'b111111100101010101111001;
         rom[873] = 24'b111111010110101111101010;
         rom[874] = 24'b111111011101110000010101;
         rom[875] = 24'b111111100001001110100111;
         rom[876] = 24'b111111101011000010101000;
         rom[877] = 24'b111111110101011100100111;
         rom[878] = 24'b111111101101101101011101;
         rom[879] = 24'b000000000100100011001110;
         rom[880] = 24'b111111110101001110000111;
         rom[881] = 24'b000000000111010010110000;
         rom[882] = 24'b000000001110001101000110;
         rom[883] = 24'b000000010010101111000111;
         rom[884] = 24'b000000010110101001001111;
         rom[885] = 24'b000000011010110100010010;
         rom[886] = 24'b000000011111100111100001;
         rom[887] = 24'b000000100000100110101011;
         rom[888] = 24'b000000011101101000110000;
         rom[889] = 24'b000000101011000011110100;
         rom[890] = 24'b000000011111001000110111;
         rom[891] = 24'b000000101010011110000101;
         rom[892] = 24'b000000100101001101110101;
         rom[893] = 24'b000000100111111111100100;
         rom[894] = 24'b000000010111001110000001;
         rom[895] = 24'b000000011111011001000010;
         rom[896] = 24'b000000001001000110111111;
         rom[897] = 24'b000000001101110000111110;
         rom[898] = 24'b000000010011111001000101;
         rom[899] = 24'b000000010011101000110100;
         rom[900] = 24'b111111111110010101001001;
         rom[901] = 24'b111111111000011110001110;
         rom[902] = 24'b111111110111111010011010;
         rom[903] = 24'b111111100111101010101100;
         rom[904] = 24'b111111011100100011001111;
         rom[905] = 24'b111111101011010111111000;
         rom[906] = 24'b111111011110001001010010;
         rom[907] = 24'b111111010101001011010100;
         rom[908] = 24'b111111011100111000001011;
         rom[909] = 24'b111111011101111000110001;
         rom[910] = 24'b111111010011101101101001;
         rom[911] = 24'b111111010010100110000010;
         rom[912] = 24'b111111100011001110011101;
         rom[913] = 24'b111111100110101011100100;
         rom[914] = 24'b111111011010111000111000;
         rom[915] = 24'b111111101110101000101000;
         rom[916] = 24'b111111101001010010100001;
         rom[917] = 24'b111111111001010100001000;
         rom[918] = 24'b111111111010100000010000;
         rom[919] = 24'b000000000000110010101111;
         rom[920] = 24'b000000000010001001001101;
         rom[921] = 24'b111111111011000000000010;
         rom[922] = 24'b000000001111010010011000;
         rom[923] = 24'b000000011001101000110101;
         rom[924] = 24'b000000010110111001011101;
         rom[925] = 24'b000000010111110110110110;
         rom[926] = 24'b000000101111001111010011;
         rom[927] = 24'b000000100000111000010110;
         rom[928] = 24'b000000100000000010011010;
         rom[929] = 24'b000000100111010100001011;
         rom[930] = 24'b000000011111001001100100;
         rom[931] = 24'b000000100111001010101100;
         rom[932] = 24'b000000011011010000111010;
         rom[933] = 24'b000000100001010001110110;
         rom[934] = 24'b000000100111100001010010;
         rom[935] = 24'b000000100001110111001011;
         rom[936] = 24'b000000010000111011010111;
         rom[937] = 24'b000000001101111010000100;
         rom[938] = 24'b000000001101101010010000;
         rom[939] = 24'b000000000111011101001010;
         rom[940] = 24'b111111111001101010000010;
         rom[941] = 24'b111111111000000101111000;
         rom[942] = 24'b111111110010001101011111;
         rom[943] = 24'b111111101100000010001100;
         rom[944] = 24'b111111101001001100001111;
         rom[945] = 24'b111111100101111001001000;
         rom[946] = 24'b111111011101000011001001;
         rom[947] = 24'b111111010111011010101100;
         rom[948] = 24'b111111011100001111000000;
         rom[949] = 24'b111111100101111010110101;
         rom[950] = 24'b111111010111001001000100;
         rom[951] = 24'b111111011000011111011011;
         rom[952] = 24'b111111010110010010001001;
         rom[953] = 24'b111111011100111001110110;
         rom[954] = 24'b111111100101111011110100;
         rom[955] = 24'b111111100100110001110101;
         rom[956] = 24'b111111101110011100101110;
         rom[957] = 24'b111111111010010010101110;
         rom[958] = 24'b111111110111101100101000;
         rom[959] = 24'b000000000001111000111010;
         rom[960] = 24'b000000001011100000101000;
         rom[961] = 24'b000000000011111001101010;
         rom[962] = 24'b000000000011101010011111;
         rom[963] = 24'b000000011011101011101110;
         rom[964] = 24'b000000011101110100001010;
         rom[965] = 24'b000000100000101111110110;
         rom[966] = 24'b000000101000001001001111;
         rom[967] = 24'b000000010101110101000111;
         rom[968] = 24'b000000011001000110000110;
         rom[969] = 24'b000000101000100110110000;
         rom[970] = 24'b000000011011000010100011;
         rom[971] = 24'b000000110000100001001000;
         rom[972] = 24'b000000101010000111011011;
         rom[973] = 24'b000000101011000001101000;
         rom[974] = 24'b000000010010100001000010;
         rom[975] = 24'b000000010111100101010000;
         rom[976] = 24'b000000011101110110010010;
         rom[977] = 24'b000000001111000101001001;
         rom[978] = 24'b000000001010100101110010;
         rom[979] = 24'b111111111100010010100101;
         rom[980] = 24'b111111111010000010100100;
         rom[981] = 24'b111111111111110111001001;
         rom[982] = 24'b111111111000011000101101;
         rom[983] = 24'b111111101100110011000111;
         rom[984] = 24'b111111101101000010110000;
         rom[985] = 24'b111111101001001111101001;
         rom[986] = 24'b111111100001101100101110;
         rom[987] = 24'b111111011101101111111110;
         rom[988] = 24'b111111010010001110001000;
         rom[989] = 24'b111111001100110101010111;
         rom[990] = 24'b111111011010101111111011;
         rom[991] = 24'b111111100001010101011001;
         rom[992] = 24'b111111010001110000000101;
         rom[993] = 24'b111111010010100101111110;
         rom[994] = 24'b111111011101010111000111;
         rom[995] = 24'b111111011111010100100000;
         rom[996] = 24'b111111110101000001101001;
         rom[997] = 24'b111111101000011110010100;
         rom[998] = 24'b000000000000011110010111;
         rom[999] = 24'b000000001001000011001010;
         rom[1000] = 24'b000000001011110100011110;
         rom[1001] = 24'b000000010010100010011110;
         rom[1002] = 24'b111111111111110010100100;
         rom[1003] = 24'b000000000100100001010111;
         rom[1004] = 24'b000000001110110010001101;
         rom[1005] = 24'b000000010001011010010100;
         rom[1006] = 24'b000000011110000000010101;
         rom[1007] = 24'b000000011111100111001110;
         rom[1008] = 24'b000000100010101110001101;
         rom[1009] = 24'b000000100111100000100100;
         rom[1010] = 24'b000000011000110110101101;
         rom[1011] = 24'b000000011111001111111100;
         rom[1012] = 24'b000000100111010111111011;
         rom[1013] = 24'b000000101000001110100111;
         rom[1014] = 24'b000000100101000000001000;
         rom[1015] = 24'b000000011111011000001111;
         rom[1016] = 24'b000000100001111110011111;
         rom[1017] = 24'b000000011100001110010001;
         rom[1018] = 24'b000000000100000001110011;
         rom[1019] = 24'b000000000100110000011011;
         rom[1020] = 24'b111111111011001011001001;
         rom[1021] = 24'b111111101101001100011000;
         rom[1022] = 24'b111111101101101000110011;
         rom[1023] = 24'b111111101001011101110111;
         rom[1024] = 24'b111111100100010011101101;
         rom[1025] = 24'b111111101010110010011111;
         rom[1026] = 24'b111111101010000101101010;
         rom[1027] = 24'b111111101101110111000011;
         rom[1028] = 24'b111111100111101100000000;
         rom[1029] = 24'b111111100001110101100010;
         rom[1030] = 24'b111111100101100001010011;
         rom[1031] = 24'b111111010011001010110100;
         rom[1032] = 24'b111111011000111001111110;
         rom[1033] = 24'b111111100001000011000000;
         rom[1034] = 24'b111111011001111011000010;
         rom[1035] = 24'b111111101101000100101001;
         rom[1036] = 24'b111111100101101100110101;
         rom[1037] = 24'b111111110110001110011100;
         rom[1038] = 24'b111111110010011000111111;
         rom[1039] = 24'b000000000001101010000111;
         rom[1040] = 24'b111111111101011100010101;
         rom[1041] = 24'b000000000111010011010111;
         rom[1042] = 24'b000000001101101001100001;
         rom[1043] = 24'b000000010111010010010101;
         rom[1044] = 24'b000000011101100010011100;
         rom[1045] = 24'b000000010111111100110001;
         rom[1046] = 24'b000000011111011100110110;
         rom[1047] = 24'b000000100011101110110101;
         rom[1048] = 24'b000000100100110011000100;
         rom[1049] = 24'b000000100101110101100000;
         rom[1050] = 24'b000000100011100001110101;
         rom[1051] = 24'b000000011111010110011101;
         rom[1052] = 24'b000000100100110001000000;
         rom[1053] = 24'b000000011101100011011101;
         rom[1054] = 24'b000000100000010011001000;
         rom[1055] = 24'b000000101000110111010011;
         rom[1056] = 24'b000000011010001111010101;
         rom[1057] = 24'b000000011010100111011000;
         rom[1058] = 24'b000000011000001000110000;
         rom[1059] = 24'b000000000001110000110011;
         rom[1060] = 24'b000000000100010011010001;
         rom[1061] = 24'b111111111010111100110101;
         rom[1062] = 24'b111111111111001000101010;
         rom[1063] = 24'b111111111001111011110111;
         rom[1064] = 24'b111111101010000101110010;
         rom[1065] = 24'b111111100110001010010111;
         rom[1066] = 24'b111111011000111101101111;
         rom[1067] = 24'b111111010111101101100100;
         rom[1068] = 24'b111111011000011110010100;
         rom[1069] = 24'b111111010111011001101110;
         rom[1070] = 24'b111111011110111011010000;
         rom[1071] = 24'b111111011001011010101000;
         rom[1072] = 24'b111111010111101011000111;
         rom[1073] = 24'b111111011101010101111010;
         rom[1074] = 24'b111111100011111010101011;
         rom[1075] = 24'b111111100110001111000000;
         rom[1076] = 24'b111111101110110111000111;
         rom[1077] = 24'b111111101111001110010000;
         rom[1078] = 24'b111111110101001011001001;
         rom[1079] = 24'b000000000100001101000001;
         rom[1080] = 24'b111111111000101101000110;
         rom[1081] = 24'b000000001101100000000011;
         rom[1082] = 24'b000000011111001110100011;
         rom[1083] = 24'b000000001011110100011100;
         rom[1084] = 24'b000000101010011010100111;
         rom[1085] = 24'b000000100001000011110010;
         rom[1086] = 24'b000000010010000010111011;
         rom[1087] = 24'b000000001100101001110011;
         rom[1088] = 24'b000000011111100100110110;
         rom[1089] = 24'b000000010111011110001110;
         rom[1090] = 24'b000000101100011000100110;
         rom[1091] = 24'b000000011101000110011000;
         rom[1092] = 24'b000000101101111110100000;
         rom[1093] = 24'b000000101100010000101001;
         rom[1094] = 24'b000000010111110101001001;
         rom[1095] = 24'b000000011000010001011100;
         rom[1096] = 24'b000000000011101100000100;
         rom[1097] = 24'b000000010101001111110110;
         rom[1098] = 24'b000000001101101001010110;
         rom[1099] = 24'b000000000010001110001101;
         rom[1100] = 24'b111111111000011010100110;
         rom[1101] = 24'b000000000001000000011101;
         rom[1102] = 24'b111111110111111011010110;
         rom[1103] = 24'b111111111000010110100110;
         rom[1104] = 24'b111111100111001111011000;
         rom[1105] = 24'b111111101001000101001010;
         rom[1106] = 24'b111111101010111100101001;
         rom[1107] = 24'b111111011001100000010010;
         rom[1108] = 24'b111111011011100011010100;
         rom[1109] = 24'b111111011010001100100000;
         rom[1110] = 24'b111111100010110100111111;
         rom[1111] = 24'b111111011010111110011001;
         rom[1112] = 24'b111111010010111100000010;
         rom[1113] = 24'b111111011001010011110011;
         rom[1114] = 24'b111111100111101101000001;
         rom[1115] = 24'b111111101110100010000101;
         rom[1116] = 24'b111111100101010010010000;
         rom[1117] = 24'b111111101111001100110010;
         rom[1118] = 24'b111111110000001001010011;
         rom[1119] = 24'b111111111101100010101001;
         rom[1120] = 24'b000000001100110011101011;
         rom[1121] = 24'b000000001111101110001011;
         rom[1122] = 24'b000000001110101000100111;
         rom[1123] = 24'b000000001001101000110001;
         rom[1124] = 24'b000000001111010010000001;
         rom[1125] = 24'b000000010101100011011101;
         rom[1126] = 24'b000000010011100100100000;
         rom[1127] = 24'b000000011101011100101011;
         rom[1128] = 24'b000000101001110101101010;
         rom[1129] = 24'b000000011001110010110110;
         rom[1130] = 24'b000000101001100010011001;
         rom[1131] = 24'b000000011110000100011110;
         rom[1132] = 24'b000000100000010010111110;
         rom[1133] = 24'b000000011100010011110100;
         rom[1134] = 24'b000000010001000010111010;
         rom[1135] = 24'b000000011100111101001001;
         rom[1136] = 24'b000000010010011011101001;
         rom[1137] = 24'b000000000010101011100011;
         rom[1138] = 24'b000000001110001101010101;
         rom[1139] = 24'b000000001011100001100011;
         rom[1140] = 24'b000000010000100011000110;
         rom[1141] = 24'b111111110101001011010111;
         rom[1142] = 24'b111111110000111101010011;
         rom[1143] = 24'b111111110000111001111010;
         rom[1144] = 24'b111111100111101010101111;
         rom[1145] = 24'b111111100111011110111001;
         rom[1146] = 24'b111111100101000001110000;
         rom[1147] = 24'b111111100000101101010110;
         rom[1148] = 24'b111111101110100101110001;
         rom[1149] = 24'b111111010011011000001000;
         rom[1150] = 24'b111111011010110001011011;
         rom[1151] = 24'b111111011101000110110101;
         rom[1152] = 24'b111111010111000110110101;
         rom[1153] = 24'b111111110000001111010001;
         rom[1154] = 24'b111111100000011001011010;
         rom[1155] = 24'b111111100000101001101001;
         rom[1156] = 24'b111111011101110101101110;
         rom[1157] = 24'b111111110010111101111010;
         rom[1158] = 24'b111111110110101000010101;
         rom[1159] = 24'b111111110110110110010010;
         rom[1160] = 24'b000000000111010010011110;
         rom[1161] = 24'b000000001110100011010001;
         rom[1162] = 24'b000000001111011001000110;
         rom[1163] = 24'b000000001010100111011000;
         rom[1164] = 24'b000000010010000110101011;
         rom[1165] = 24'b000000010111001010100010;
         rom[1166] = 24'b000000101000000010101010;
         rom[1167] = 24'b000000101010110111110011;
         rom[1168] = 24'b000000101100011001110101;
         rom[1169] = 24'b000000110000010000101100;
         rom[1170] = 24'b000000011100111000110011;
         rom[1171] = 24'b000000100100000011110000;
         rom[1172] = 24'b000000010110111000010111;
         rom[1173] = 24'b000000101011110110000011;
         rom[1174] = 24'b000000011100001001111010;
         rom[1175] = 24'b000000011010101010001101;
         rom[1176] = 24'b000000011011101000011111;
         rom[1177] = 24'b000000001011100110000111;
         rom[1178] = 24'b000000001010010110100100;
         rom[1179] = 24'b000000000101111110011101;
         rom[1180] = 24'b000000000001011110110100;
         rom[1181] = 24'b111111111001100011111101;
         rom[1182] = 24'b111111110110101010101101;
         rom[1183] = 24'b111111101110111011110101;
         rom[1184] = 24'b111111101011010111100100;
         rom[1185] = 24'b111111101011000001000011;
         rom[1186] = 24'b111111100001011011101110;
         rom[1187] = 24'b111111010110110101000000;
         rom[1188] = 24'b111111011110100100000100;
         rom[1189] = 24'b111111011100101011101111;
         rom[1190] = 24'b111111010010111111100011;
         rom[1191] = 24'b111111011000111011000010;
         rom[1192] = 24'b111111100100001110110001;
         rom[1193] = 24'b111111011001001011111101;
         rom[1194] = 24'b111111100000110110011000;
         rom[1195] = 24'b111111100010001101010010;
         rom[1196] = 24'b111111100000111100110101;
         rom[1197] = 24'b111111100101011001001100;
         rom[1198] = 24'b111111110100011001010010;
         rom[1199] = 24'b111111111000110101000011;
         rom[1200] = 24'b111111111101101010010011;
         rom[1201] = 24'b000000001110010111011101;
         rom[1202] = 24'b000000010000111101100011;
         rom[1203] = 24'b000000011010101101010110;
         rom[1204] = 24'b000000011101100100000011;
         rom[1205] = 24'b000000100001010100001011;
         rom[1206] = 24'b000000011010011111001101;
         rom[1207] = 24'b000000011111000111111100;
         rom[1208] = 24'b000000011001000010100000;
         rom[1209] = 24'b000000100101010011000001;
         rom[1210] = 24'b000000011110110100111001;
         rom[1211] = 24'b000000100110011000110111;
         rom[1212] = 24'b000000100011101101111100;
         rom[1213] = 24'b000000110000100011100001;
         rom[1214] = 24'b000000100101010100001111;
         rom[1215] = 24'b000000010111101011011111;
         rom[1216] = 24'b000000001100010111000101;
         rom[1217] = 24'b000000000011101000010000;
         rom[1218] = 24'b000000001101100001100100;
         rom[1219] = 24'b000000001110000010110000;
         rom[1220] = 24'b111111111111111001111111;
         rom[1221] = 24'b111111110011000001111010;
         rom[1222] = 24'b111111101000000011000110;
         rom[1223] = 24'b111111100111011101001000;
         rom[1224] = 24'b111111101100100000101111;
         rom[1225] = 24'b111111100100101111011110;
         rom[1226] = 24'b111111100000011110001001;
         rom[1227] = 24'b111111101110100010111000;
         rom[1228] = 24'b111111100100000100101011;
         rom[1229] = 24'b111111100010001001010000;
         rom[1230] = 24'b111111010111000011010011;
         rom[1231] = 24'b111111101000001011110101;
         rom[1232] = 24'b111111101010111110111010;
         rom[1233] = 24'b111111100000011111100101;
         rom[1234] = 24'b111111100101100010011010;
         rom[1235] = 24'b111111100000111110011011;
         rom[1236] = 24'b111111101001111101101011;
         rom[1237] = 24'b111111110101011010000111;
         rom[1238] = 24'b111111110100101011110110;
         rom[1239] = 24'b111111111011000101000100;
         rom[1240] = 24'b000000001011101000001101;
         rom[1241] = 24'b000000000000010101011100;
         rom[1242] = 24'b000000000101111110001111;
         rom[1243] = 24'b000000011100100001110011;
         rom[1244] = 24'b000000010101110000011110;
         rom[1245] = 24'b000000010111101010111001;
         rom[1246] = 24'b000000010111000000100010;
         rom[1247] = 24'b000000101001000111001111;
         rom[1248] = 24'b000000100101011110001110;
         rom[1249] = 24'b000000100100101011110101;
         rom[1250] = 24'b000000100001010000001011;
         rom[1251] = 24'b000000011110011010010010;
         rom[1252] = 24'b000000011101110101100100;
         rom[1253] = 24'b000000100010110000000111;
         rom[1254] = 24'b000000100001001011110001;
         rom[1255] = 24'b000000010011001100010000;
         rom[1256] = 24'b000000010110000100111101;
         rom[1257] = 24'b000000000100111100101000;
         rom[1258] = 24'b000000000110111110011100;
         rom[1259] = 24'b000000000010001111011101;
         rom[1260] = 24'b111111110111000011111010;
         rom[1261] = 24'b111111111011100101001101;
         rom[1262] = 24'b111111101111001011010110;
         rom[1263] = 24'b111111101010100010111010;
         rom[1264] = 24'b111111100110111010110011;
         rom[1265] = 24'b111111100101010010000110;
         rom[1266] = 24'b111111011110011100101000;
         rom[1267] = 24'b111111100000111100011100;
         rom[1268] = 24'b111111010011111100010011;
         rom[1269] = 24'b111111101010101111001001;
         rom[1270] = 24'b111111100000100101111011;
         rom[1271] = 24'b111111001111010010110110;
         rom[1272] = 24'b111111011011000101010001;
         rom[1273] = 24'b111111011101100011000110;
         rom[1274] = 24'b111111101011111011010011;
         rom[1275] = 24'b111111100111011100000110;
         rom[1276] = 24'b111111101111100101001100;
         rom[1277] = 24'b111111101010000101001100;
         rom[1278] = 24'b111111110101100110010101;
         rom[1279] = 24'b111111111001101001110110;
         rom[1280] = 24'b111111111111010111110101;
         rom[1281] = 24'b000000001010111011010010;
         rom[1282] = 24'b000000000001110011010000;
         rom[1283] = 24'b000000010000010110110111;
         rom[1284] = 24'b000000101000001100001101;
         rom[1285] = 24'b000000010111101010001111;
         rom[1286] = 24'b000000100111111110101001;
         rom[1287] = 24'b000000100001000111010110;
         rom[1288] = 24'b000000011001111000100001;
         rom[1289] = 24'b000000100000101000111000;
         rom[1290] = 24'b000000100101111110011001;
         rom[1291] = 24'b000000011110110110010100;
         rom[1292] = 24'b000000100100111101111000;
         rom[1293] = 24'b000000101001100001010011;
         rom[1294] = 24'b000000100011101001011001;
         rom[1295] = 24'b000000010000110011101100;
         rom[1296] = 24'b000000011001110001000101;
         rom[1297] = 24'b000000011100101111010010;
         rom[1298] = 24'b000000010000100100000110;
         rom[1299] = 24'b000000001000100100111000;
         rom[1300] = 24'b111111110011111010001111;
         rom[1301] = 24'b111111111011011000000011;
         rom[1302] = 24'b000000001000010110001100;
         rom[1303] = 24'b000000001000111011111010;
         rom[1304] = 24'b000000000110000111111000;
         rom[1305] = 24'b000000001100001110100000;
         rom[1306] = 24'b000000001000111111110000;
         rom[1307] = 24'b000000010100111011111001;
         rom[1308] = 24'b000000001100111101100001;
         rom[1309] = 24'b000000100001001100001000;
         rom[1310] = 24'b000000100111101001110101;
         rom[1311] = 24'b000000101001100100001010;
         rom[1312] = 24'b000000111100001110011100;
         rom[1313] = 24'b000000110110100111111111;
         rom[1314] = 24'b000001001011000011001110;
         rom[1315] = 24'b000001010110101011110101;
         rom[1316] = 24'b000001100100000011010110;
         rom[1317] = 24'b000001110101110100001000;
         rom[1318] = 24'b000001111100110111111100;
         rom[1319] = 24'b000010001010001100011101;
         rom[1320] = 24'b000010010100001011111101;
         rom[1321] = 24'b000010010111011011010101;
         rom[1322] = 24'b000010101100100110100001;
         rom[1323] = 24'b000010110011110111101010;
         rom[1324] = 24'b000011000100110110010001;
         rom[1325] = 24'b000011010101011011000100;
         rom[1326] = 24'b000011010101100011101010;
         rom[1327] = 24'b000011100011110001010010;
         rom[1328] = 24'b000011100101010010101111;
         rom[1329] = 24'b000100000001001000001000;
         rom[1330] = 24'b000100000111010101111100;
         rom[1331] = 24'b000100000110010110111101;
         rom[1332] = 24'b000100001000000010001100;
         rom[1333] = 24'b000100001100011100101000;
         rom[1334] = 24'b000100010110010111101111;
         rom[1335] = 24'b000100010110111011110111;
         rom[1336] = 24'b000100001011011011000100;
         rom[1337] = 24'b000100100111010111111010;
         rom[1338] = 24'b000100011111100101001010;
         rom[1339] = 24'b000100011100000010011100;
         rom[1340] = 24'b000100101010000010110111;
         rom[1341] = 24'b000100100100101001101111;
         rom[1342] = 24'b000100011100110100101011;
         rom[1343] = 24'b000100100101101110101101;
         rom[1344] = 24'b000100101100101110101100;
         rom[1345] = 24'b000100101000110011100010;
         rom[1346] = 24'b000100111010111010100111;
         rom[1347] = 24'b000100110111001111000101;
         rom[1348] = 24'b000100111001001010110101;
         rom[1349] = 24'b000100111111011111110000;
         rom[1350] = 24'b000101010100111000000110;
         rom[1351] = 24'b000101000100010001100010;
         rom[1352] = 24'b000101011011001001000010;
         rom[1353] = 24'b000101110010111001011100;
         rom[1354] = 24'b000101100100000010010100;
         rom[1355] = 24'b000101111010110101001111;
         rom[1356] = 24'b000101111101010110010100;
         rom[1357] = 24'b000110001101000110100011;
         rom[1358] = 24'b000110011000110000100000;
         rom[1359] = 24'b000110100001101011111110;
         rom[1360] = 24'b000110101110001111101101;
         rom[1361] = 24'b000111001010011101101011;
         rom[1362] = 24'b000111010110100111010100;
         rom[1363] = 24'b000111011110111001010101;
         rom[1364] = 24'b000111101000101010100111;
         rom[1365] = 24'b000111101111100101000010;
         rom[1366] = 24'b000111110110001100011000;
         rom[1367] = 24'b001000000001001111111100;
         rom[1368] = 24'b001000100010011010101101;
         rom[1369] = 24'b001000011010010011111010;
         rom[1370] = 24'b001000100110111010111110;
         rom[1371] = 24'b001000101000000000001101;
         rom[1372] = 24'b001000101011110110101001;
         rom[1373] = 24'b001000111110101110001111;
         rom[1374] = 24'b001000110101010010111011;
         rom[1375] = 24'b001001001100000110110110;
         rom[1376] = 24'b001000111010101010100001;
         rom[1377] = 24'b001000110011011011000100;
         rom[1378] = 24'b001000111111010010010001;
         rom[1379] = 24'b001000111110011101001101;
         rom[1380] = 24'b001001001110000000001110;
         rom[1381] = 24'b001001001011001001111101;
         rom[1382] = 24'b001001000100100100111100;
         rom[1383] = 24'b001001001100011001100101;
         rom[1384] = 24'b001001010000110011101100;
         rom[1385] = 24'b001001001111101000001101;
         rom[1386] = 24'b001001011010011001100010;
         rom[1387] = 24'b001001011011111111000110;
         rom[1388] = 24'b001001011010110000011001;
         rom[1389] = 24'b001001001100100000101100;
         rom[1390] = 24'b001001001100100101111110;
         rom[1391] = 24'b001000110110001001111011;
         rom[1392] = 24'b001000111000111001001111;
         rom[1393] = 24'b001000101101100011000101;
         rom[1394] = 24'b001000101101000101111101;
         rom[1395] = 24'b001000110101010011111111;
         rom[1396] = 24'b001000101100001010010000;
         rom[1397] = 24'b001000101111100111111101;
         rom[1398] = 24'b001000101000101100001110;
         rom[1399] = 24'b001000011111001000011001;
         rom[1400] = 24'b001000100010100001010011;
         rom[1401] = 24'b001000010110010011111111;
         rom[1402] = 24'b001000010011010111010011;
         rom[1403] = 24'b001000101111000111010111;
         rom[1404] = 24'b001000010101110001011111;
         rom[1405] = 24'b001000011010011000101110;
         rom[1406] = 24'b001000001011111010010101;
         rom[1407] = 24'b001000010111010111111000;
         rom[1408] = 24'b001000010000010010100000;
         rom[1409] = 24'b001000001100000110110110;
         rom[1410] = 24'b001000000000000111010000;
         rom[1411] = 24'b000111101111001110001011;
         rom[1412] = 24'b000111111110100101000000;
         rom[1413] = 24'b000111010111110100101011;
         rom[1414] = 24'b000111010101010100011010;
         rom[1415] = 24'b000111010110011100011011;
         rom[1416] = 24'b000111000010110110010011;
         rom[1417] = 24'b000110111110001000110111;
         rom[1418] = 24'b000110110001010100110011;
         rom[1419] = 24'b000110011001001010100010;
         rom[1420] = 24'b000110011000110101101101;
         rom[1421] = 24'b000110000010111101010110;
         rom[1422] = 24'b000101110000010010100101;
         rom[1423] = 24'b000101110010100001000111;
         rom[1424] = 24'b000101100111100000011101;
         rom[1425] = 24'b000101011000001101101010;
         rom[1426] = 24'b000101001000011010010100;
         rom[1427] = 24'b000100110101000111000101;
         rom[1428] = 24'b000100111000111011111001;
         rom[1429] = 24'b000100101111011101100010;
         rom[1430] = 24'b000100100010101101000101;
         rom[1431] = 24'b000100011100001111011101;
         rom[1432] = 24'b000100011011011010010100;
         rom[1433] = 24'b000100001111110101011101;
         rom[1434] = 24'b000100010001100001000000;
         rom[1435] = 24'b000100001011001111011000;
         rom[1436] = 24'b000100001010100110110111;
         rom[1437] = 24'b000100000110110010100110;
         rom[1438] = 24'b000100000110011011111110;
         rom[1439] = 24'b000100000100011011111100;
         rom[1440] = 24'b000100001000111010100101;
         rom[1441] = 24'b000100001010010000010100;
         rom[1442] = 24'b000100000100010111011101;
         rom[1443] = 24'b000011110110001101100000;
         rom[1444] = 24'b000011110110101011111000;
         rom[1445] = 24'b000011101111110010110000;
         rom[1446] = 24'b000011110111110100111110;
         rom[1447] = 24'b000011101110010000101111;
         rom[1448] = 24'b000011110001011110001110;
         rom[1449] = 24'b000011011011111110100011;
         rom[1450] = 24'b000011100010000101011111;
         rom[1451] = 24'b000011011000001010001110;
         rom[1452] = 24'b000010111110100111000101;
         rom[1453] = 24'b000011010000011100011101;
         rom[1454] = 24'b000010111011111010110110;
         rom[1455] = 24'b000010110000101100101110;
         rom[1456] = 24'b000010100001010101011001;
         rom[1457] = 24'b000010010110101000001101;
         rom[1458] = 24'b000010001001010111010000;
         rom[1459] = 24'b000001110010111111100110;
         rom[1460] = 24'b000001100101110000100100;
         rom[1461] = 24'b000001011100111111001111;
         rom[1462] = 24'b000001100110100100110110;
         rom[1463] = 24'b000001001101001001101101;
         rom[1464] = 24'b000001000001110101101000;
         rom[1465] = 24'b000000101110111011010100;
         rom[1466] = 24'b000000101100101011010010;
         rom[1467] = 24'b000000011111101000010011;
         rom[1468] = 24'b000000001001111010110011;
         rom[1469] = 24'b000000001101010110111101;
         rom[1470] = 24'b000000000110110011010100;
         rom[1471] = 24'b111111101111011110110110;
         rom[1472] = 24'b111111110111010101100100;
         rom[1473] = 24'b111111100010100001101101;
         rom[1474] = 24'b111111100111000100100001;
         rom[1475] = 24'b111111100000011001011100;
         rom[1476] = 24'b111111100100110111101111;
         rom[1477] = 24'b111111101010000010101011;
         rom[1478] = 24'b111111100110010100111111;
         rom[1479] = 24'b111111100101110000101001;
         rom[1480] = 24'b111111011001010000111011;
         rom[1481] = 24'b111111010101101011011100;
         rom[1482] = 24'b111111100100001100010011;
         rom[1483] = 24'b111111011011100101101100;
         rom[1484] = 24'b111111010101100110111010;
         rom[1485] = 24'b111111010110011101100011;
         rom[1486] = 24'b111110111111110010010010;
         rom[1487] = 24'b111111001010101100010101;
         rom[1488] = 24'b111111001101010111000100;
         rom[1489] = 24'b111111011001011011100111;
         rom[1490] = 24'b111111010110000111010001;
         rom[1491] = 24'b111111011111011010100101;
         rom[1492] = 24'b111111110000100101000010;
         rom[1493] = 24'b111111101110111100110101;
         rom[1494] = 24'b111111101110000101111110;
         rom[1495] = 24'b111111111001011111001011;
         rom[1496] = 24'b111111101011000101001000;
         rom[1497] = 24'b111111111001100001001101;
         rom[1498] = 24'b111111111100001111111111;
         rom[1499] = 24'b111111111100001110110010;
         rom[1500] = 24'b111111111110000101001010;
         rom[1501] = 24'b111111111000010011011111;
         rom[1502] = 24'b111111111011011110101010;
         rom[1503] = 24'b111111110011011010000101;
         rom[1504] = 24'b111111101111110110111000;
         rom[1505] = 24'b111111101000111111010010;
         rom[1506] = 24'b111111011010001001111110;
         rom[1507] = 24'b111111101011010001000011;
         rom[1508] = 24'b111111001101100110001110;
         rom[1509] = 24'b111111100010011110100000;
         rom[1510] = 24'b111111011101010111111111;
         rom[1511] = 24'b111111010100111011100100;
         rom[1512] = 24'b111111011110110110111111;
         rom[1513] = 24'b111111100110010100000010;
         rom[1514] = 24'b111111011100100110010111;
         rom[1515] = 24'b111111101010001100000101;
         rom[1516] = 24'b111111101000100100110001;
         rom[1517] = 24'b111111101001110101001101;
         rom[1518] = 24'b111111111000110111111101;
         rom[1519] = 24'b111111111101100001000001;
         rom[1520] = 24'b000000000000111001100110;
         rom[1521] = 24'b000000001100011010010101;
         rom[1522] = 24'b000000010011100010110010;
         rom[1523] = 24'b000000010000000101010000;
         rom[1524] = 24'b000000010000110001111101;
         rom[1525] = 24'b000000011100101101011000;
         rom[1526] = 24'b000000011010011100110110;
         rom[1527] = 24'b000000011011010001100101;
         rom[1528] = 24'b000000100100001111101111;
         rom[1529] = 24'b000000011100011110000110;
         rom[1530] = 24'b000000110011001101111111;
         rom[1531] = 24'b000000101101110001100011;
         rom[1532] = 24'b000000100100001111101110;
         rom[1533] = 24'b000000100000110101111110;
         rom[1534] = 24'b000000011100001000011101;
         rom[1535] = 24'b000000100010001001011100;
         rom[1536] = 24'b000000010110010011000001;
         rom[1537] = 24'b000000001011011100100100;
         rom[1538] = 24'b000000001000100111000101;
         rom[1539] = 24'b000000001010110101011001;
         rom[1540] = 24'b000000000111101101100110;
         rom[1541] = 24'b111111111001010100111000;
         rom[1542] = 24'b111111110001110110001110;
         rom[1543] = 24'b111111101101100100101100;
         rom[1544] = 24'b111111110011100110111111;
         rom[1545] = 24'b111111011000001011010000;
         rom[1546] = 24'b111111100010011100111001;
         rom[1547] = 24'b111111100101001010011101;
         rom[1548] = 24'b111111001101111100000111;
         rom[1549] = 24'b111111011111011101111111;
         rom[1550] = 24'b111111100001100000100000;
         rom[1551] = 24'b111111001010011111011010;
         rom[1552] = 24'b111111010111111011000001;
         rom[1553] = 24'b111111011010000010001111;
         rom[1554] = 24'b111111010110001010110011;
         rom[1555] = 24'b111111100110000110010101;
         rom[1556] = 24'b111111101111010000010110;
         rom[1557] = 24'b111111111000110011100100;
         rom[1558] = 24'b000000000111001011011001;
         rom[1559] = 24'b000000000111001110100101;
         rom[1560] = 24'b111111111010111101010001;
         rom[1561] = 24'b000000000000101010110001;
         rom[1562] = 24'b000000001111000110101000;
         rom[1563] = 24'b000000010001001001001111;
         rom[1564] = 24'b000000011011111100000110;
         rom[1565] = 24'b000000010111101000000011;
         rom[1566] = 24'b000000011001000110010100;
         rom[1567] = 24'b000000100010111110010111;
         rom[1568] = 24'b000000010111001000010101;
         rom[1569] = 24'b000000100011110111000010;
         rom[1570] = 24'b000000101010110100101110;
         rom[1571] = 24'b000000101011111010000010;
         rom[1572] = 24'b000000011110100000010011;
         rom[1573] = 24'b000000100011111001101111;
         rom[1574] = 24'b000000100001001000110000;
         rom[1575] = 24'b000000011010001111110101;
         rom[1576] = 24'b000000001110101101000101;
         rom[1577] = 24'b000000000110011110110111;
         rom[1578] = 24'b000000000001111100100100;
         rom[1579] = 24'b000000001001010000101001;
         rom[1580] = 24'b000000001000010110100000;
         rom[1581] = 24'b000000000000010011011011;
         rom[1582] = 24'b111111110111011010001000;
         rom[1583] = 24'b111111100111100000101010;
         rom[1584] = 24'b111111100111100101111111;
         rom[1585] = 24'b111111100101011000010000;
         rom[1586] = 24'b111111011000111011000000;
         rom[1587] = 24'b111111100001110101100010;
         rom[1588] = 24'b111111100101000100101001;
         rom[1589] = 24'b111111010000100101100010;
         rom[1590] = 24'b111111011010100011110000;
         rom[1591] = 24'b111111011111100011101011;
         rom[1592] = 24'b111111011001101100001101;
         rom[1593] = 24'b111111011101101000111001;
         rom[1594] = 24'b111111101101010000000111;
         rom[1595] = 24'b111111100100111110001110;
         rom[1596] = 24'b111111101010100001011000;
         rom[1597] = 24'b000000000100000000111010;
         rom[1598] = 24'b111111101010101000011011;
         rom[1599] = 24'b111111110100110100100111;
         rom[1600] = 24'b111111110110111000011101;
         rom[1601] = 24'b000000000011110001111000;
         rom[1602] = 24'b000000010100111010111010;
         rom[1603] = 24'b000000001111000101001101;
         rom[1604] = 24'b000000010101000011000001;
         rom[1605] = 24'b000000011110010111100000;
         rom[1606] = 24'b000000011011111010101101;
         rom[1607] = 24'b000000101000110101010110;
         rom[1608] = 24'b000000100101010111100101;
         rom[1609] = 24'b000000100010011000111010;
         rom[1610] = 24'b000000011100100111110110;
         rom[1611] = 24'b000000100001001000111000;
         rom[1612] = 24'b000000011000101101000011;
         rom[1613] = 24'b000000011001100000100101;
         rom[1614] = 24'b000000010010001100110110;
         rom[1615] = 24'b000000011000100010010101;
         rom[1616] = 24'b000000010100100011011000;
         rom[1617] = 24'b000000001100000010011100;
         rom[1618] = 24'b000000000101111010111101;
         rom[1619] = 24'b000000001010110001010101;
         rom[1620] = 24'b111111111110100011110101;
         rom[1621] = 24'b000000000100100111111011;
         rom[1622] = 24'b111111110101101111001111;
         rom[1623] = 24'b111111111100010100111110;
         rom[1624] = 24'b111111101110100011001010;
         rom[1625] = 24'b111111101010110011000101;
         rom[1626] = 24'b111111100101010101010100;
         rom[1627] = 24'b111111101100010001001010;
         rom[1628] = 24'b111111101001110000100110;
         rom[1629] = 24'b111111011101101110110001;
         rom[1630] = 24'b111111011010011010000011;
         rom[1631] = 24'b111111011000100001101110;
         rom[1632] = 24'b111111101000101010101010;
         rom[1633] = 24'b111111101100011011011101;
         rom[1634] = 24'b111111011101011010001010;
         rom[1635] = 24'b111111010011110000010111;
         rom[1636] = 24'b111111100010000111010001;
         rom[1637] = 24'b111111111011010010110110;
         rom[1638] = 24'b111111110000110111110100;
         rom[1639] = 24'b111111111100000100001001;
         rom[1640] = 24'b111111111110001011001110;
         rom[1641] = 24'b000000010001010011001010;
         rom[1642] = 24'b000000011100110111000010;
         rom[1643] = 24'b000000010111000111000000;
         rom[1644] = 24'b000000101101000000111010;
         rom[1645] = 24'b000000111110011100111010;
         rom[1646] = 24'b000000111100100000000111;
         rom[1647] = 24'b000001000000110011101000;
         rom[1648] = 24'b000000110011111100100001;
         rom[1649] = 24'b000001001001011000011001;
         rom[1650] = 24'b000001001111000010100111;
         rom[1651] = 24'b000001010100110000010100;
         rom[1652] = 24'b000001010010100000100100;
         rom[1653] = 24'b000001001011111100010001;
         rom[1654] = 24'b000001010010110000101001;
         rom[1655] = 24'b000001000110001101111110;
         rom[1656] = 24'b000001001001010101011010;
         rom[1657] = 24'b000000111100010101001010;
         rom[1658] = 24'b000000111000111010011011;
         rom[1659] = 24'b000001000000010111000010;
         rom[1660] = 24'b000000110000101100001110;
         rom[1661] = 24'b000000110111011101001000;
         rom[1662] = 24'b000000100110100000000011;
         rom[1663] = 24'b000000100101111111111000;
         rom[1664] = 24'b000000101001011100111000;
         rom[1665] = 24'b000000010011100001100101;
         rom[1666] = 24'b000000011100000101101000;
         rom[1667] = 24'b000000101010101001010100;
         rom[1668] = 24'b000000010100011010011011;
         rom[1669] = 24'b000000110001000001010111;
         rom[1670] = 24'b000000011011111000010001;
         rom[1671] = 24'b000000011101000111011111;
         rom[1672] = 24'b000000011100010011001111;
         rom[1673] = 24'b000000011101010110101000;
         rom[1674] = 24'b000000101001001101010000;
         rom[1675] = 24'b000000101101100000101001;
         rom[1676] = 24'b000000111010100010111100;
         rom[1677] = 24'b000000110110011111101111;
         rom[1678] = 24'b000000111110111110001110;
         rom[1679] = 24'b000000111100100011100000;
         rom[1680] = 24'b000001001101000111010000;
         rom[1681] = 24'b000001011111011110101100;
         rom[1682] = 24'b000001010101001010001001;
         rom[1683] = 24'b000001001110110010111110;
         rom[1684] = 24'b000001100001000011010001;
         rom[1685] = 24'b000001010111101111001101;
         rom[1686] = 24'b000001100011111011100011;
         rom[1687] = 24'b000001111001101111110010;
         rom[1688] = 24'b000001101010101100011011;
         rom[1689] = 24'b000001111010101000111011;
         rom[1690] = 24'b000001111100111110001110;
         rom[1691] = 24'b000010000000001011010000;
         rom[1692] = 24'b000001111010101000100111;
         rom[1693] = 24'b000001101111010000010111;
         rom[1694] = 24'b000001111001001100000000;
         rom[1695] = 24'b000001110101000101110100;
         rom[1696] = 24'b000001110000011101101100;
         rom[1697] = 24'b000001101100001011000100;
         rom[1698] = 24'b000001100001101010011010;
         rom[1699] = 24'b000001100110001100011000;
         rom[1700] = 24'b000001011001110010000111;
         rom[1701] = 24'b000001100000111010101100;
         rom[1702] = 24'b000001010010001000110111;
         rom[1703] = 24'b000001001010010111100101;
         rom[1704] = 24'b000001001111011010000110;
         rom[1705] = 24'b000000111101001000001110;
         rom[1706] = 24'b000001000010111100111110;
         rom[1707] = 24'b000000111111111100000111;
         rom[1708] = 24'b000000111001011000111100;
         rom[1709] = 24'b000001000111110000101110;
         rom[1710] = 24'b000001000100011011110111;
         rom[1711] = 24'b000001000110001110000010;
         rom[1712] = 24'b000000110111101010101110;
         rom[1713] = 24'b000001001000000001100011;
         rom[1714] = 24'b000001001011111011000011;
         rom[1715] = 24'b000001011010100001101101;
         rom[1716] = 24'b000001010000110101111010;
         rom[1717] = 24'b000001001110010101110111;
         rom[1718] = 24'b000001010010010000001100;
         rom[1719] = 24'b000001011101001111101101;
         rom[1720] = 24'b000001100100101101100111;
         rom[1721] = 24'b000001101100111011010000;
         rom[1722] = 24'b000001110101001111111000;
         rom[1723] = 24'b000001110011111001101010;
         rom[1724] = 24'b000001111000011101011110;
         rom[1725] = 24'b000010000000000011110001;
         rom[1726] = 24'b000001111100100111101111;
         rom[1727] = 24'b000001111111010100001000;
         rom[1728] = 24'b000010010101110011001110;
         rom[1729] = 24'b000010001101100011001111;
         rom[1730] = 24'b000010010111111111110001;
         rom[1731] = 24'b000010001100100010100111;
         rom[1732] = 24'b000010001110101001011101;
         rom[1733] = 24'b000010001100111010111110;
         rom[1734] = 24'b000010000011111011011100;
         rom[1735] = 24'b000010010010111100010011;
         rom[1736] = 24'b000001111110100100000110;
         rom[1737] = 24'b000001110110010111101101;
         rom[1738] = 24'b000001110001100110011111;
         rom[1739] = 24'b000001101100111000000110;
         rom[1740] = 24'b000001100101010101011110;
         rom[1741] = 24'b000001101111100100111111;
         rom[1742] = 24'b000001100001110000111100;
         rom[1743] = 24'b000001101111101110111011;
         rom[1744] = 24'b000001011000000010011010;
         rom[1745] = 24'b000001100001001011010011;
         rom[1746] = 24'b000001001100000111101000;
         rom[1747] = 24'b000001010001001000111100;
         rom[1748] = 24'b000001000111010110000010;
         rom[1749] = 24'b000001000110011001000110;
         rom[1750] = 24'b000001000110010011010101;
         rom[1751] = 24'b000001001100001111010011;
         rom[1752] = 24'b000001010011110011101010;
         rom[1753] = 24'b000001001110010000010111;
         rom[1754] = 24'b000001000100000010111000;
         rom[1755] = 24'b000001001010111010100000;
         rom[1756] = 24'b000001011011111010011011;
         rom[1757] = 24'b000001010101100011011011;
         rom[1758] = 24'b000001101110110100001001;
         rom[1759] = 24'b000001111100011001010010;
         rom[1760] = 24'b000001101011111011010101;
         rom[1761] = 24'b000010000110110010001000;
         rom[1762] = 24'b000010000000010101111111;
         rom[1763] = 24'b000001111011110000101110;
         rom[1764] = 24'b000001111110001001000010;
         rom[1765] = 24'b000010010000101000011010;
         rom[1766] = 24'b000010001000001110100101;
         rom[1767] = 24'b000010010000101100100011;
         rom[1768] = 24'b000010011010101001100100;
         rom[1769] = 24'b000010011001111000101000;
         rom[1770] = 24'b000010011010001000001110;
         rom[1771] = 24'b000010100010000001011110;
         rom[1772] = 24'b000010011110110110010101;
         rom[1773] = 24'b000010001100001111001001;
         rom[1774] = 24'b000010011101100000110110;
         rom[1775] = 24'b000010010001110100100101;
         rom[1776] = 24'b000010001101011000100010;
         rom[1777] = 24'b000010001101011000011010;
         rom[1778] = 24'b000001111100111011010111;
         rom[1779] = 24'b000001110110111101110100;
         rom[1780] = 24'b000010000110000010111001;
         rom[1781] = 24'b000001110100110010010000;
         rom[1782] = 24'b000001100111000011101000;
         rom[1783] = 24'b000001011101010110001000;
         rom[1784] = 24'b000001110010111110000101;
         rom[1785] = 24'b000001011011110100010111;
         rom[1786] = 24'b000001011000011010111000;
         rom[1787] = 24'b000001001011000001000010;
         rom[1788] = 24'b000001001110100110011011;
         rom[1789] = 24'b000001010000000110111000;
         rom[1790] = 24'b000001011111100110100110;
         rom[1791] = 24'b000001010000110101101001;
         rom[1792] = 24'b000001010110111000110100;
         rom[1793] = 24'b000001010111000001110101;
         rom[1794] = 24'b000001010101000011100100;
         rom[1795] = 24'b000001011110000000100000;
         rom[1796] = 24'b000001011110000011100010;
         rom[1797] = 24'b000001101110011100001110;
         rom[1798] = 24'b000001100101000010100110;
         rom[1799] = 24'b000001101011011010100100;
         rom[1800] = 24'b000001110101001001110111;
         rom[1801] = 24'b000001111100100010110110;
         rom[1802] = 24'b000001111110111000011100;
         rom[1803] = 24'b000010001010000111100000;
         rom[1804] = 24'b000010001111000111100011;
         rom[1805] = 24'b000010001101101011100000;
         rom[1806] = 24'b000010001111000011011010;
         rom[1807] = 24'b000010100111111110011100;
         rom[1808] = 24'b000010100110000101011111;
         rom[1809] = 24'b000010100000001000111000;
         rom[1810] = 24'b000010010110011000011001;
         rom[1811] = 24'b000010011111000101110111;
         rom[1812] = 24'b000010101000111100000001;
         rom[1813] = 24'b000010001110010101111010;
         rom[1814] = 24'b000010001111100101101111;
         rom[1815] = 24'b000010010000111010001011;
         rom[1816] = 24'b000010010101010011101000;
         rom[1817] = 24'b000010001010001010100100;
         rom[1818] = 24'b000001111001000011010100;
         rom[1819] = 24'b000010001000001100000111;
         rom[1820] = 24'b000001100101110110011001;
         rom[1821] = 24'b000001111011011001110001;
         rom[1822] = 24'b000001111001110001011110;
         rom[1823] = 24'b000001101110110100001101;
         rom[1824] = 24'b000001011110000001001110;
         rom[1825] = 24'b000001100011100000010100;
         rom[1826] = 24'b000001100011001000010101;
         rom[1827] = 24'b000001001011101110110100;
         rom[1828] = 24'b000001000101110100101100;
         rom[1829] = 24'b000001011110011111100001;
         rom[1830] = 24'b000001001010011011111111;
         rom[1831] = 24'b000001010110001110000101;
         rom[1832] = 24'b000001010010011110001100;
         rom[1833] = 24'b000001011000111110111010;
         rom[1834] = 24'b000001010001010100110111;
         rom[1835] = 24'b000001011100001011011111;
         rom[1836] = 24'b000001100100010101011110;
         rom[1837] = 24'b000001100111011100000111;
         rom[1838] = 24'b000001110100011000111110;
         rom[1839] = 24'b000010000000111001001000;
         rom[1840] = 24'b000001110101111011101011;
         rom[1841] = 24'b000010000000101011111010;
         rom[1842] = 24'b000010000011111100101001;
         rom[1843] = 24'b000010000111001110110111;
         rom[1844] = 24'b000010010010011111010010;
         rom[1845] = 24'b000010001000011100010010;
         rom[1846] = 24'b000010100010011000010101;
         rom[1847] = 24'b000010011011111101010101;
         rom[1848] = 24'b000010001100111000001110;
         rom[1849] = 24'b000010011011001001111000;
         rom[1850] = 24'b000010011111101010101000;
         rom[1851] = 24'b000010010100010111011000;
         rom[1852] = 24'b000010101010110101010111;
         rom[1853] = 24'b000010010010100001111101;
         rom[1854] = 24'b000010001011001111001101;
         rom[1855] = 24'b000010010101110011001001;
         rom[1856] = 24'b000010000111100110110001;
         rom[1857] = 24'b000010001000011111001010;
         rom[1858] = 24'b000010000011111011100010;
         rom[1859] = 24'b000010000011011011110111;
         rom[1860] = 24'b000001110100001000111011;
         rom[1861] = 24'b000001110111000011100110;
         rom[1862] = 24'b000001100101011110101000;
         rom[1863] = 24'b000001011111000001100101;
         rom[1864] = 24'b000001100101001000010111;
         rom[1865] = 24'b000001011100000100000011;
         rom[1866] = 24'b000001010000011000110101;
         rom[1867] = 24'b000001011001110001101001;
         rom[1868] = 24'b000001011100011101100111;
         rom[1869] = 24'b000001010011011101111111;
         rom[1870] = 24'b000001010011000110010110;
         rom[1871] = 24'b000001000110001100110010;
         rom[1872] = 24'b000001011000111101101110;
         rom[1873] = 24'b000001010111011110101110;
         rom[1874] = 24'b000001011101100011100101;
         rom[1875] = 24'b000001001110001011110011;
         rom[1876] = 24'b000001101011100001111010;
         rom[1877] = 24'b000001110011111111111101;
         rom[1878] = 24'b000001101011010111001110;
         rom[1879] = 24'b000001111110100011101101;
         rom[1880] = 24'b000001111011001100001101;
         rom[1881] = 24'b000001111110000110100010;
         rom[1882] = 24'b000001111000110111000111;
         rom[1883] = 24'b000010001000100011101000;
         rom[1884] = 24'b000010010011111000110101;
         rom[1885] = 24'b000010000111010101110101;
         rom[1886] = 24'b000010001101101100001101;
         rom[1887] = 24'b000010011011111100010010;
         rom[1888] = 24'b000010010111110001111110;
         rom[1889] = 24'b000010001110000011011011;
         rom[1890] = 24'b000010100100011001001001;
         rom[1891] = 24'b000010001100111101011000;
         rom[1892] = 24'b000010010100111100001011;
         rom[1893] = 24'b000010000101011010011000;
         rom[1894] = 24'b000010010011000100111110;
         rom[1895] = 24'b000010010000001111011001;
         rom[1896] = 24'b000001111010101100011110;
         rom[1897] = 24'b000001110001001100010001;
         rom[1898] = 24'b000001110010011101000101;
         rom[1899] = 24'b000001110100000100001111;
         rom[1900] = 24'b000001101010000001011000;
         rom[1901] = 24'b000001100001101100010111;
         rom[1902] = 24'b000001101000011010111011;
         rom[1903] = 24'b000001100001000101110101;
         rom[1904] = 24'b000001000101101010010001;
         rom[1905] = 24'b000001011010000010011010;
         rom[1906] = 24'b000001010001000011100001;
         rom[1907] = 24'b000001010111001100111100;
         rom[1908] = 24'b000000111110010001001101;
         rom[1909] = 24'b000001000011001000010010;
         rom[1910] = 24'b000000111110111110111110;
         rom[1911] = 24'b000001001001001001111001;
         rom[1912] = 24'b000000111110001011101010;
         rom[1913] = 24'b000001001110001111000100;
         rom[1914] = 24'b000001000100010101001111;
         rom[1915] = 24'b000001010001000010010001;
         rom[1916] = 24'b000001001110010000101000;
         rom[1917] = 24'b000001001111010100000100;
         rom[1918] = 24'b000001001100010001101100;
         rom[1919] = 24'b000001011101000110000100;
         rom[1920] = 24'b000001100011010110001001;
         rom[1921] = 24'b000001101101111000001011;
         rom[1922] = 24'b000001100010101011001100;
         rom[1923] = 24'b000001111001011101100101;
         rom[1924] = 24'b000010000010001101001010;
         rom[1925] = 24'b000010000100111100101101;
         rom[1926] = 24'b000010000101101110110100;
         rom[1927] = 24'b000010000000101011000000;
         rom[1928] = 24'b000001110011000101010111;
         rom[1929] = 24'b000010000110000111101000;
         rom[1930] = 24'b000010001100000100100101;
         rom[1931] = 24'b000010000110111110101011;
         rom[1932] = 24'b000010000011110001000111;
         rom[1933] = 24'b000001110111010100000101;
         rom[1934] = 24'b000010000100000010010101;
         rom[1935] = 24'b000010000100001100000000;
         rom[1936] = 24'b000001111110111001110101;
         rom[1937] = 24'b000001101001111001110001;
         rom[1938] = 24'b000001110000100001000001;
         rom[1939] = 24'b000001011110000010001111;
         rom[1940] = 24'b000001011000111101010010;
         rom[1941] = 24'b000001010001100011111110;
         rom[1942] = 24'b000001001000101110010010;
         rom[1943] = 24'b000001001110011111001101;
         rom[1944] = 24'b000001010000100110001100;
         rom[1945] = 24'b000000110110010001110001;
         rom[1946] = 24'b000000101110011001110101;
         rom[1947] = 24'b000000110100101001101110;
         rom[1948] = 24'b000000110110010001011011;
         rom[1949] = 24'b000000101110000100001110;
         rom[1950] = 24'b000000101110010101000011;
         rom[1951] = 24'b000001000000001101000110;
         rom[1952] = 24'b000000101110001110111010;
         rom[1953] = 24'b000000101101101010001100;
         rom[1954] = 24'b000000110011010110000011;
         rom[1955] = 24'b000000110100110000011110;
         rom[1956] = 24'b000000101101101100110100;
         rom[1957] = 24'b000001000010110100111110;
         rom[1958] = 24'b000001000111000101011011;
         rom[1959] = 24'b000001010110111010110101;
         rom[1960] = 24'b000001000101100101010101;
         rom[1961] = 24'b000001010011000100011101;
         rom[1962] = 24'b000001010011101010100001;
         rom[1963] = 24'b000001011111110010110100;
         rom[1964] = 24'b000001100010110110111010;
         rom[1965] = 24'b000001001100110001011101;
         rom[1966] = 24'b000001011100100100000101;
         rom[1967] = 24'b000001101001011111100001;
         rom[1968] = 24'b000001101000001000110010;
         rom[1969] = 24'b000001101001010011001100;
         rom[1970] = 24'b000001101100011100101111;
         rom[1971] = 24'b000001101111111000101011;
         rom[1972] = 24'b000001011000100000000010;
         rom[1973] = 24'b000001100001011100100101;
         rom[1974] = 24'b000001100100001000110010;
         rom[1975] = 24'b000001100001100101110111;
         rom[1976] = 24'b000001011010111101011101;
         rom[1977] = 24'b000001010101010111000100;
         rom[1978] = 24'b000000111111111011100110;
         rom[1979] = 24'b000000111001111101110011;
         rom[1980] = 24'b000000110110000000011111;
         rom[1981] = 24'b000000101111010110111110;
         rom[1982] = 24'b000000100101010101000110;
         rom[1983] = 24'b000000100000101101010110;
         rom[1984] = 24'b000000011110001010100011;
         rom[1985] = 24'b000000011011011010111100;
         rom[1986] = 24'b000000011011101101011001;
         rom[1987] = 24'b000000001011100010111000;
         rom[1988] = 24'b111111111001000110100000;
         rom[1989] = 24'b111111111011100011110100;
         rom[1990] = 24'b111111110100010100010111;
         rom[1991] = 24'b000000001100100111010101;
         rom[1992] = 24'b111111110111011000010110;
         rom[1993] = 24'b000000001110110000011101;
         rom[1994] = 24'b111111111000000111010110;
         rom[1995] = 24'b000000001010010110101110;
         rom[1996] = 24'b111111111101111110001101;
         rom[1997] = 24'b000000010010001000111001;
         rom[1998] = 24'b000000000001000100111110;
         rom[1999] = 24'b000000000010011010010010;
         end 

	 always @(posedge(clk))
		 begin 
			 if(reset) 
				 begin 
					 data_out <= 24'b0; 
					 i <= 16'b0; 
					 counter <= 16'b0; 
				 end 
			 else 
				 begin 
					 if(counter == 16'd5000) 
						 begin 
							 data_out <= rom[i]; 
							 counter <=16'b0; 
							 if(i == 1999) i <= 0; 
							 else i <= i + 1; 
						 end 
					 else counter <= counter + 16'd1; 
				 end 
		 end 

endmodule
