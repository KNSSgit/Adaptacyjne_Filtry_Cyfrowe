`timescale 1ns/100ps

module gen_sinus( 
 	 output reg signed [23:0] data_out,
	 input clk,
	 input reset
	 ); 

	 reg signed [23:0] rom[0:959];
	 reg [15:0] i;
	 reg [15:0] counter;

	 always @(reset)
		 begin 
			 rom[0] = 24'b000000000000000000000000;
			 rom[1] = 24'b001010101011100110000000;
			 rom[2] = 24'b010010100000000001001110;
			 rom[3] = 24'b010101010111001100000000;
			 rom[4] = 24'b010010100000000001001110;
			 rom[5] = 24'b001010101011100110000000;
			 rom[6] = 24'b000000000000000000000000;
			 rom[7] = 24'b110101010100011010000000;
			 rom[8] = 24'b101101011111111110110010;
			 rom[9] = 24'b101010101000110100000000;
			 rom[10] = 24'b101101011111111110110010;
			 rom[11] = 24'b110101010100011010000000;
			 rom[12] = 24'b000000000000000000000000;
			 rom[13] = 24'b001010101011100110000000;
			 rom[14] = 24'b010010100000000001001110;
			 rom[15] = 24'b010101010111001100000000;
			 rom[16] = 24'b010010100000000001001110;
			 rom[17] = 24'b001010101011100110000000;
			 rom[18] = 24'b000000000000000000000000;
			 rom[19] = 24'b110101010100011010000000;
			 rom[20] = 24'b101101011111111110110010;
			 rom[21] = 24'b101010101000110100000000;
			 rom[22] = 24'b101101011111111110110010;
			 rom[23] = 24'b110101010100011010000000;
			 rom[24] = 24'b000000000000000000000000;
			 rom[25] = 24'b001010101011100110000000;
			 rom[26] = 24'b010010100000000001001110;
			 rom[27] = 24'b010101010111001100000000;
			 rom[28] = 24'b010010100000000001001110;
			 rom[29] = 24'b001010101011100110000000;
			 rom[30] = 24'b000000000000000000000000;
			 rom[31] = 24'b110101010100011010000000;
			 rom[32] = 24'b101101011111111110110010;
			 rom[33] = 24'b101010101000110100000000;
			 rom[34] = 24'b101101011111111110110010;
			 rom[35] = 24'b110101010100011010000000;
			 rom[36] = 24'b000000000000000000000000;
			 rom[37] = 24'b001010101011100110000000;
			 rom[38] = 24'b010010100000000001001110;
			 rom[39] = 24'b010101010111001100000000;
			 rom[40] = 24'b010010100000000001001110;
			 rom[41] = 24'b001010101011100110000000;
			 rom[42] = 24'b000000000000000000000000;
			 rom[43] = 24'b110101010100011010000000;
			 rom[44] = 24'b101101011111111110110010;
			 rom[45] = 24'b101010101000110100000000;
			 rom[46] = 24'b101101011111111110110010;
			 rom[47] = 24'b110101010100011010000000;
			 rom[48] = 24'b000000000000000000000000;
			 rom[49] = 24'b001010101011100110000000;
			 rom[50] = 24'b010010100000000001001110;
			 rom[51] = 24'b010101010111001100000000;
			 rom[52] = 24'b010010100000000001001110;
			 rom[53] = 24'b001010101011100110000000;
			 rom[54] = 24'b000000000000000000000000;
			 rom[55] = 24'b110101010100011010000000;
			 rom[56] = 24'b101101011111111110110010;
			 rom[57] = 24'b101010101000110100000000;
			 rom[58] = 24'b101101011111111110110010;
			 rom[59] = 24'b110101010100011010000000;
			 rom[60] = 24'b000000000000000000000000;
			 rom[61] = 24'b001010101011100110000000;
			 rom[62] = 24'b010010100000000001001110;
			 rom[63] = 24'b010101010111001100000000;
			 rom[64] = 24'b010010100000000001001110;
			 rom[65] = 24'b001010101011100110000000;
			 rom[66] = 24'b000000000000000000000000;
			 rom[67] = 24'b110101010100011010000000;
			 rom[68] = 24'b101101011111111110110010;
			 rom[69] = 24'b101010101000110100000000;
			 rom[70] = 24'b101101011111111110110010;
			 rom[71] = 24'b110101010100011010000000;
			 rom[72] = 24'b000000000000000000000000;
			 rom[73] = 24'b001010101011100110000000;
			 rom[74] = 24'b010010100000000001001110;
			 rom[75] = 24'b010101010111001100000000;
			 rom[76] = 24'b010010100000000001001110;
			 rom[77] = 24'b001010101011100110000000;
			 rom[78] = 24'b000000000000000000000000;
			 rom[79] = 24'b110101010100011010000000;
			 rom[80] = 24'b101101011111111110110010;
			 rom[81] = 24'b101010101000110100000000;
			 rom[82] = 24'b101101011111111110110010;
			 rom[83] = 24'b110101010100011010000000;
			 rom[84] = 24'b000000000000000000000000;
			 rom[85] = 24'b001010101011100110000000;
			 rom[86] = 24'b010010100000000001001110;
			 rom[87] = 24'b010101010111001100000000;
			 rom[88] = 24'b010010100000000001001110;
			 rom[89] = 24'b001010101011100110000000;
			 rom[90] = 24'b000000000000000000000000;
			 rom[91] = 24'b110101010100011010000000;
			 rom[92] = 24'b101101011111111110110010;
			 rom[93] = 24'b101010101000110100000000;
			 rom[94] = 24'b101101011111111110110010;
			 rom[95] = 24'b110101010100011010000000;
			 rom[96] = 24'b000000000000000000000000;
			 rom[97] = 24'b001010101011100110000000;
			 rom[98] = 24'b010010100000000001001110;
			 rom[99] = 24'b010101010111001100000000;
			 rom[100] = 24'b010010100000000001001110;
			 rom[101] = 24'b001010101011100110000000;
			 rom[102] = 24'b000000000000000000000000;
			 rom[103] = 24'b110101010100011010000000;
			 rom[104] = 24'b101101011111111110110010;
			 rom[105] = 24'b101010101000110100000000;
			 rom[106] = 24'b101101011111111110110010;
			 rom[107] = 24'b110101010100011010000000;
			 rom[108] = 24'b000000000000000000000000;
			 rom[109] = 24'b001010101011100110000000;
			 rom[110] = 24'b010010100000000001001110;
			 rom[111] = 24'b010101010111001100000000;
			 rom[112] = 24'b010010100000000001001110;
			 rom[113] = 24'b001010101011100110000000;
			 rom[114] = 24'b000000000000000000000000;
			 rom[115] = 24'b110101010100011010000000;
			 rom[116] = 24'b101101011111111110110010;
			 rom[117] = 24'b101010101000110100000000;
			 rom[118] = 24'b101101011111111110110010;
			 rom[119] = 24'b110101010100011010000000;
			 rom[120] = 24'b000000000000000000000000;
			 rom[121] = 24'b001010101011100110000000;
			 rom[122] = 24'b010010100000000001001110;
			 rom[123] = 24'b010101010111001100000000;
			 rom[124] = 24'b010010100000000001001110;
			 rom[125] = 24'b001010101011100110000000;
			 rom[126] = 24'b000000000000000000000000;
			 rom[127] = 24'b110101010100011010000000;
			 rom[128] = 24'b101101011111111110110010;
			 rom[129] = 24'b101010101000110100000000;
			 rom[130] = 24'b101101011111111110110010;
			 rom[131] = 24'b110101010100011010000000;
			 rom[132] = 24'b000000000000000000000000;
			 rom[133] = 24'b001010101011100110000000;
			 rom[134] = 24'b010010100000000001001110;
			 rom[135] = 24'b010101010111001100000000;
			 rom[136] = 24'b010010100000000001001110;
			 rom[137] = 24'b001010101011100110000000;
			 rom[138] = 24'b000000000000000000000000;
			 rom[139] = 24'b110101010100011010000000;
			 rom[140] = 24'b101101011111111110110010;
			 rom[141] = 24'b101010101000110100000000;
			 rom[142] = 24'b101101011111111110110010;
			 rom[143] = 24'b110101010100011010000000;
			 rom[144] = 24'b000000000000000000000000;
			 rom[145] = 24'b001010101011100110000000;
			 rom[146] = 24'b010010100000000001001110;
			 rom[147] = 24'b010101010111001100000000;
			 rom[148] = 24'b010010100000000001001110;
			 rom[149] = 24'b001010101011100110000000;
			 rom[150] = 24'b000000000000000000000000;
			 rom[151] = 24'b110101010100011010000000;
			 rom[152] = 24'b101101011111111110110010;
			 rom[153] = 24'b101010101000110100000000;
			 rom[154] = 24'b101101011111111110110010;
			 rom[155] = 24'b110101010100011010000000;
			 rom[156] = 24'b000000000000000000000000;
			 rom[157] = 24'b001010101011100110000000;
			 rom[158] = 24'b010010100000000001001110;
			 rom[159] = 24'b010101010111001100000000;
			 rom[160] = 24'b010010100000000001001110;
			 rom[161] = 24'b001010101011100110000000;
			 rom[162] = 24'b000000000000000000000000;
			 rom[163] = 24'b110101010100011010000000;
			 rom[164] = 24'b101101011111111110110010;
			 rom[165] = 24'b101010101000110100000000;
			 rom[166] = 24'b101101011111111110110010;
			 rom[167] = 24'b110101010100011010000000;
			 rom[168] = 24'b000000000000000000000000;
			 rom[169] = 24'b001010101011100110000000;
			 rom[170] = 24'b010010100000000001001110;
			 rom[171] = 24'b010101010111001100000000;
			 rom[172] = 24'b010010100000000001001110;
			 rom[173] = 24'b001010101011100110000000;
			 rom[174] = 24'b000000000000000000000000;
			 rom[175] = 24'b110101010100011010000000;
			 rom[176] = 24'b101101011111111110110010;
			 rom[177] = 24'b101010101000110100000000;
			 rom[178] = 24'b101101011111111110110010;
			 rom[179] = 24'b110101010100011010000000;
			 rom[180] = 24'b000000000000000000000000;
			 rom[181] = 24'b001010101011100110000000;
			 rom[182] = 24'b010010100000000001001110;
			 rom[183] = 24'b010101010111001100000000;
			 rom[184] = 24'b010010100000000001001110;
			 rom[185] = 24'b001010101011100110000000;
			 rom[186] = 24'b000000000000000000000000;
			 rom[187] = 24'b110101010100011010000000;
			 rom[188] = 24'b101101011111111110110010;
			 rom[189] = 24'b101010101000110100000000;
			 rom[190] = 24'b101101011111111110110010;
			 rom[191] = 24'b110101010100011010000000;
			 rom[192] = 24'b000000000000000000000000;
			 rom[193] = 24'b001010101011100110000000;
			 rom[194] = 24'b010010100000000001001110;
			 rom[195] = 24'b010101010111001100000000;
			 rom[196] = 24'b010010100000000001001110;
			 rom[197] = 24'b001010101011100110000000;
			 rom[198] = 24'b000000000000000000000000;
			 rom[199] = 24'b110101010100011010000000;
			 rom[200] = 24'b101101011111111110110010;
			 rom[201] = 24'b101010101000110100000000;
			 rom[202] = 24'b101101011111111110110010;
			 rom[203] = 24'b110101010100011010000000;
			 rom[204] = 24'b000000000000000000000000;
			 rom[205] = 24'b001010101011100110000000;
			 rom[206] = 24'b010010100000000001001110;
			 rom[207] = 24'b010101010111001100000000;
			 rom[208] = 24'b010010100000000001001110;
			 rom[209] = 24'b001010101011100110000000;
			 rom[210] = 24'b000000000000000000000000;
			 rom[211] = 24'b110101010100011010000000;
			 rom[212] = 24'b101101011111111110110010;
			 rom[213] = 24'b101010101000110100000000;
			 rom[214] = 24'b101101011111111110110010;
			 rom[215] = 24'b110101010100011010000000;
			 rom[216] = 24'b000000000000000000000000;
			 rom[217] = 24'b001010101011100110000000;
			 rom[218] = 24'b010010100000000001001110;
			 rom[219] = 24'b010101010111001100000000;
			 rom[220] = 24'b010010100000000001001110;
			 rom[221] = 24'b001010101011100110000000;
			 rom[222] = 24'b000000000000000000000000;
			 rom[223] = 24'b110101010100011010000000;
			 rom[224] = 24'b101101011111111110110010;
			 rom[225] = 24'b101010101000110100000000;
			 rom[226] = 24'b101101011111111110110010;
			 rom[227] = 24'b110101010100011010000000;
			 rom[228] = 24'b000000000000000000000000;
			 rom[229] = 24'b001010101011100110000000;
			 rom[230] = 24'b010010100000000001001110;
			 rom[231] = 24'b010101010111001100000000;
			 rom[232] = 24'b010010100000000001001110;
			 rom[233] = 24'b001010101011100110000000;
			 rom[234] = 24'b000000000000000000000000;
			 rom[235] = 24'b110101010100011010000000;
			 rom[236] = 24'b101101011111111110110010;
			 rom[237] = 24'b101010101000110100000000;
			 rom[238] = 24'b101101011111111110110010;
			 rom[239] = 24'b110101010100011010000000;
			 rom[240] = 24'b000000000000000000000000;
			 rom[241] = 24'b001010101011100110000000;
			 rom[242] = 24'b010010100000000001001110;
			 rom[243] = 24'b010101010111001100000000;
			 rom[244] = 24'b010010100000000001001110;
			 rom[245] = 24'b001010101011100110000000;
			 rom[246] = 24'b000000000000000000000000;
			 rom[247] = 24'b110101010100011010000000;
			 rom[248] = 24'b101101011111111110110010;
			 rom[249] = 24'b101010101000110100000000;
			 rom[250] = 24'b101101011111111110110010;
			 rom[251] = 24'b110101010100011010000000;
			 rom[252] = 24'b000000000000000000000000;
			 rom[253] = 24'b001010101011100110000000;
			 rom[254] = 24'b010010100000000001001110;
			 rom[255] = 24'b010101010111001100000000;
			 rom[256] = 24'b010010100000000001001110;
			 rom[257] = 24'b001010101011100110000000;
			 rom[258] = 24'b000000000000000000000000;
			 rom[259] = 24'b110101010100011010000000;
			 rom[260] = 24'b101101011111111110110010;
			 rom[261] = 24'b101010101000110100000000;
			 rom[262] = 24'b101101011111111110110010;
			 rom[263] = 24'b110101010100011010000000;
			 rom[264] = 24'b000000000000000000000000;
			 rom[265] = 24'b001010101011100110000000;
			 rom[266] = 24'b010010100000000001001110;
			 rom[267] = 24'b010101010111001100000000;
			 rom[268] = 24'b010010100000000001001110;
			 rom[269] = 24'b001010101011100110000000;
			 rom[270] = 24'b000000000000000000000000;
			 rom[271] = 24'b110101010100011010000000;
			 rom[272] = 24'b101101011111111110110010;
			 rom[273] = 24'b101010101000110100000000;
			 rom[274] = 24'b101101011111111110110010;
			 rom[275] = 24'b110101010100011010000000;
			 rom[276] = 24'b000000000000000000000000;
			 rom[277] = 24'b001010101011100110000000;
			 rom[278] = 24'b010010100000000001001110;
			 rom[279] = 24'b010101010111001100000000;
			 rom[280] = 24'b010010100000000001001110;
			 rom[281] = 24'b001010101011100110000000;
			 rom[282] = 24'b000000000000000000000000;
			 rom[283] = 24'b110101010100011010000000;
			 rom[284] = 24'b101101011111111110110010;
			 rom[285] = 24'b101010101000110100000000;
			 rom[286] = 24'b101101011111111110110010;
			 rom[287] = 24'b110101010100011010000000;
			 rom[288] = 24'b000000000000000000000000;
			 rom[289] = 24'b001010101011100110000000;
			 rom[290] = 24'b010010100000000001001110;
			 rom[291] = 24'b010101010111001100000000;
			 rom[292] = 24'b010010100000000001001110;
			 rom[293] = 24'b001010101011100110000000;
			 rom[294] = 24'b000000000000000000000000;
			 rom[295] = 24'b110101010100011010000000;
			 rom[296] = 24'b101101011111111110110010;
			 rom[297] = 24'b101010101000110100000000;
			 rom[298] = 24'b101101011111111110110010;
			 rom[299] = 24'b110101010100011010000000;
			 rom[300] = 24'b000000000000000000000000;
			 rom[301] = 24'b001010101011100110000000;
			 rom[302] = 24'b010010100000000001001110;
			 rom[303] = 24'b010101010111001100000000;
			 rom[304] = 24'b010010100000000001001110;
			 rom[305] = 24'b001010101011100110000000;
			 rom[306] = 24'b000000000000000000000000;
			 rom[307] = 24'b110101010100011010000000;
			 rom[308] = 24'b101101011111111110110010;
			 rom[309] = 24'b101010101000110100000000;
			 rom[310] = 24'b101101011111111110110010;
			 rom[311] = 24'b110101010100011010000000;
			 rom[312] = 24'b000000000000000000000000;
			 rom[313] = 24'b001010101011100110000000;
			 rom[314] = 24'b010010100000000001001110;
			 rom[315] = 24'b010101010111001100000000;
			 rom[316] = 24'b010010100000000001001110;
			 rom[317] = 24'b001010101011100110000000;
			 rom[318] = 24'b000000000000000000000000;
			 rom[319] = 24'b110101010100011010000000;
			 rom[320] = 24'b101101011111111110110010;
			 rom[321] = 24'b101010101000110100000000;
			 rom[322] = 24'b101101011111111110110010;
			 rom[323] = 24'b110101010100011010000000;
			 rom[324] = 24'b000000000000000000000000;
			 rom[325] = 24'b001010101011100110000000;
			 rom[326] = 24'b010010100000000001001110;
			 rom[327] = 24'b010101010111001100000000;
			 rom[328] = 24'b010010100000000001001110;
			 rom[329] = 24'b001010101011100110000000;
			 rom[330] = 24'b000000000000000000000000;
			 rom[331] = 24'b110101010100011010000000;
			 rom[332] = 24'b101101011111111110110010;
			 rom[333] = 24'b101010101000110100000000;
			 rom[334] = 24'b101101011111111110110010;
			 rom[335] = 24'b110101010100011010000000;
			 rom[336] = 24'b000000000000000000000000;
			 rom[337] = 24'b001010101011100110000000;
			 rom[338] = 24'b010010100000000001001110;
			 rom[339] = 24'b010101010111001100000000;
			 rom[340] = 24'b010010100000000001001110;
			 rom[341] = 24'b001010101011100110000000;
			 rom[342] = 24'b000000000000000000000000;
			 rom[343] = 24'b110101010100011010000000;
			 rom[344] = 24'b101101011111111110110010;
			 rom[345] = 24'b101010101000110100000000;
			 rom[346] = 24'b101101011111111110110010;
			 rom[347] = 24'b110101010100011010000000;
			 rom[348] = 24'b000000000000000000000000;
			 rom[349] = 24'b001010101011100110000000;
			 rom[350] = 24'b010010100000000001001110;
			 rom[351] = 24'b010101010111001100000000;
			 rom[352] = 24'b010010100000000001001110;
			 rom[353] = 24'b001010101011100110000000;
			 rom[354] = 24'b000000000000000000000000;
			 rom[355] = 24'b110101010100011010000000;
			 rom[356] = 24'b101101011111111110110010;
			 rom[357] = 24'b101010101000110100000000;
			 rom[358] = 24'b101101011111111110110010;
			 rom[359] = 24'b110101010100011010000000;
			 rom[360] = 24'b000000000000000000000000;
			 rom[361] = 24'b001010101011100110000000;
			 rom[362] = 24'b010010100000000001001110;
			 rom[363] = 24'b010101010111001100000000;
			 rom[364] = 24'b010010100000000001001110;
			 rom[365] = 24'b001010101011100110000000;
			 rom[366] = 24'b000000000000000000000000;
			 rom[367] = 24'b110101010100011010000000;
			 rom[368] = 24'b101101011111111110110010;
			 rom[369] = 24'b101010101000110100000000;
			 rom[370] = 24'b101101011111111110110010;
			 rom[371] = 24'b110101010100011010000000;
			 rom[372] = 24'b000000000000000000000000;
			 rom[373] = 24'b001010101011100110000000;
			 rom[374] = 24'b010010100000000001001110;
			 rom[375] = 24'b010101010111001100000000;
			 rom[376] = 24'b010010100000000001001110;
			 rom[377] = 24'b001010101011100110000000;
			 rom[378] = 24'b000000000000000000000000;
			 rom[379] = 24'b110101010100011010000000;
			 rom[380] = 24'b101101011111111110110010;
			 rom[381] = 24'b101010101000110100000000;
			 rom[382] = 24'b101101011111111110110010;
			 rom[383] = 24'b110101010100011010000000;
			 rom[384] = 24'b000000000000000000000000;
			 rom[385] = 24'b001010101011100110000000;
			 rom[386] = 24'b010010100000000001001110;
			 rom[387] = 24'b010101010111001100000000;
			 rom[388] = 24'b010010100000000001001110;
			 rom[389] = 24'b001010101011100110000000;
			 rom[390] = 24'b000000000000000000000000;
			 rom[391] = 24'b110101010100011010000000;
			 rom[392] = 24'b101101011111111110110010;
			 rom[393] = 24'b101010101000110100000000;
			 rom[394] = 24'b101101011111111110110010;
			 rom[395] = 24'b110101010100011010000000;
			 rom[396] = 24'b000000000000000000000000;
			 rom[397] = 24'b001010101011100110000000;
			 rom[398] = 24'b010010100000000001001110;
			 rom[399] = 24'b010101010111001100000000;
			 rom[400] = 24'b010010100000000001001110;
			 rom[401] = 24'b001010101011100110000000;
			 rom[402] = 24'b000000000000000000000000;
			 rom[403] = 24'b110101010100011010000000;
			 rom[404] = 24'b101101011111111110110010;
			 rom[405] = 24'b101010101000110100000000;
			 rom[406] = 24'b101101011111111110110010;
			 rom[407] = 24'b110101010100011010000000;
			 rom[408] = 24'b000000000000000000000000;
			 rom[409] = 24'b001010101011100110000000;
			 rom[410] = 24'b010010100000000001001110;
			 rom[411] = 24'b010101010111001100000000;
			 rom[412] = 24'b010010100000000001001110;
			 rom[413] = 24'b001010101011100110000000;
			 rom[414] = 24'b000000000000000000000000;
			 rom[415] = 24'b110101010100011010000000;
			 rom[416] = 24'b101101011111111110110010;
			 rom[417] = 24'b101010101000110100000000;
			 rom[418] = 24'b101101011111111110110010;
			 rom[419] = 24'b110101010100011010000000;
			 rom[420] = 24'b000000000000000000000000;
			 rom[421] = 24'b001010101011100110000000;
			 rom[422] = 24'b010010100000000001001110;
			 rom[423] = 24'b010101010111001100000000;
			 rom[424] = 24'b010010100000000001001110;
			 rom[425] = 24'b001010101011100110000000;
			 rom[426] = 24'b000000000000000000000000;
			 rom[427] = 24'b110101010100011010000000;
			 rom[428] = 24'b101101011111111110110010;
			 rom[429] = 24'b101010101000110100000000;
			 rom[430] = 24'b101101011111111110110010;
			 rom[431] = 24'b110101010100011010000000;
			 rom[432] = 24'b000000000000000000000000;
			 rom[433] = 24'b001010101011100110000000;
			 rom[434] = 24'b010010100000000001001110;
			 rom[435] = 24'b010101010111001100000000;
			 rom[436] = 24'b010010100000000001001110;
			 rom[437] = 24'b001010101011100110000000;
			 rom[438] = 24'b000000000000000000000000;
			 rom[439] = 24'b110101010100011010000000;
			 rom[440] = 24'b101101011111111110110010;
			 rom[441] = 24'b101010101000110100000000;
			 rom[442] = 24'b101101011111111110110010;
			 rom[443] = 24'b110101010100011010000000;
			 rom[444] = 24'b000000000000000000000000;
			 rom[445] = 24'b001010101011100110000000;
			 rom[446] = 24'b010010100000000001001110;
			 rom[447] = 24'b010101010111001100000000;
			 rom[448] = 24'b010010100000000001001110;
			 rom[449] = 24'b001010101011100110000000;
			 rom[450] = 24'b000000000000000000000000;
			 rom[451] = 24'b110101010100011010000000;
			 rom[452] = 24'b101101011111111110110010;
			 rom[453] = 24'b101010101000110100000000;
			 rom[454] = 24'b101101011111111110110010;
			 rom[455] = 24'b110101010100011010000000;
			 rom[456] = 24'b000000000000000000000000;
			 rom[457] = 24'b001010101011100110000000;
			 rom[458] = 24'b010010100000000001001110;
			 rom[459] = 24'b010101010111001100000000;
			 rom[460] = 24'b010010100000000001001110;
			 rom[461] = 24'b001010101011100110000000;
			 rom[462] = 24'b000000000000000000000000;
			 rom[463] = 24'b110101010100011010000000;
			 rom[464] = 24'b101101011111111110110010;
			 rom[465] = 24'b101010101000110100000000;
			 rom[466] = 24'b101101011111111110110010;
			 rom[467] = 24'b110101010100011010000000;
			 rom[468] = 24'b000000000000000000000000;
			 rom[469] = 24'b001010101011100110000000;
			 rom[470] = 24'b010010100000000001001110;
			 rom[471] = 24'b010101010111001100000000;
			 rom[472] = 24'b010010100000000001001110;
			 rom[473] = 24'b001010101011100110000000;
			 rom[474] = 24'b000000000000000000000000;
			 rom[475] = 24'b110101010100011010000000;
			 rom[476] = 24'b101101011111111110110010;
			 rom[477] = 24'b101010101000110100000000;
			 rom[478] = 24'b101101011111111110110010;
			 rom[479] = 24'b110101010100011010000000;
			 rom[480] = 24'b000000000000000000000000;
			 rom[481] = 24'b001010101011100110000000;
			 rom[482] = 24'b010010100000000001001110;
			 rom[483] = 24'b010101010111001100000000;
			 rom[484] = 24'b010010100000000001001110;
			 rom[485] = 24'b001010101011100110000000;
			 rom[486] = 24'b000000000000000000000000;
			 rom[487] = 24'b110101010100011010000000;
			 rom[488] = 24'b101101011111111110110010;
			 rom[489] = 24'b101010101000110100000000;
			 rom[490] = 24'b101101011111111110110010;
			 rom[491] = 24'b110101010100011010000000;
			 rom[492] = 24'b000000000000000000000000;
			 rom[493] = 24'b001010101011100110000000;
			 rom[494] = 24'b010010100000000001001110;
			 rom[495] = 24'b010101010111001100000000;
			 rom[496] = 24'b010010100000000001001110;
			 rom[497] = 24'b001010101011100110000000;
			 rom[498] = 24'b000000000000000000000000;
			 rom[499] = 24'b110101010100011010000000;
			 rom[500] = 24'b101101011111111110110010;
			 rom[501] = 24'b101010101000110100000000;
			 rom[502] = 24'b101101011111111110110010;
			 rom[503] = 24'b110101010100011010000000;
			 rom[504] = 24'b000000000000000000000000;
			 rom[505] = 24'b001010101011100110000000;
			 rom[506] = 24'b010010100000000001001110;
			 rom[507] = 24'b010101010111001100000000;
			 rom[508] = 24'b010010100000000001001110;
			 rom[509] = 24'b001010101011100110000000;
			 rom[510] = 24'b000000000000000000000000;
			 rom[511] = 24'b110101010100011010000000;
			 rom[512] = 24'b101101011111111110110010;
			 rom[513] = 24'b101010101000110100000000;
			 rom[514] = 24'b101101011111111110110010;
			 rom[515] = 24'b110101010100011010000000;
			 rom[516] = 24'b000000000000000000000000;
			 rom[517] = 24'b001010101011100110000000;
			 rom[518] = 24'b010010100000000001001110;
			 rom[519] = 24'b010101010111001100000000;
			 rom[520] = 24'b010010100000000001001110;
			 rom[521] = 24'b001010101011100110000000;
			 rom[522] = 24'b000000000000000000000000;
			 rom[523] = 24'b110101010100011010000000;
			 rom[524] = 24'b101101011111111110110010;
			 rom[525] = 24'b101010101000110100000000;
			 rom[526] = 24'b101101011111111110110010;
			 rom[527] = 24'b110101010100011010000000;
			 rom[528] = 24'b000000000000000000000000;
			 rom[529] = 24'b001010101011100110000000;
			 rom[530] = 24'b010010100000000001001110;
			 rom[531] = 24'b010101010111001100000000;
			 rom[532] = 24'b010010100000000001001110;
			 rom[533] = 24'b001010101011100110000000;
			 rom[534] = 24'b000000000000000000000000;
			 rom[535] = 24'b110101010100011010000000;
			 rom[536] = 24'b101101011111111110110010;
			 rom[537] = 24'b101010101000110100000000;
			 rom[538] = 24'b101101011111111110110010;
			 rom[539] = 24'b110101010100011010000000;
			 rom[540] = 24'b000000000000000000000000;
			 rom[541] = 24'b001010101011100110000000;
			 rom[542] = 24'b010010100000000001001110;
			 rom[543] = 24'b010101010111001100000000;
			 rom[544] = 24'b010010100000000001001110;
			 rom[545] = 24'b001010101011100110000000;
			 rom[546] = 24'b000000000000000000000000;
			 rom[547] = 24'b110101010100011010000000;
			 rom[548] = 24'b101101011111111110110010;
			 rom[549] = 24'b101010101000110100000000;
			 rom[550] = 24'b101101011111111110110010;
			 rom[551] = 24'b110101010100011010000000;
			 rom[552] = 24'b000000000000000000000000;
			 rom[553] = 24'b001010101011100110000000;
			 rom[554] = 24'b010010100000000001001110;
			 rom[555] = 24'b010101010111001100000000;
			 rom[556] = 24'b010010100000000001001110;
			 rom[557] = 24'b001010101011100110000000;
			 rom[558] = 24'b000000000000000000000000;
			 rom[559] = 24'b110101010100011010000000;
			 rom[560] = 24'b101101011111111110110010;
			 rom[561] = 24'b101010101000110100000000;
			 rom[562] = 24'b101101011111111110110010;
			 rom[563] = 24'b110101010100011010000000;
			 rom[564] = 24'b000000000000000000000000;
			 rom[565] = 24'b001010101011100110000000;
			 rom[566] = 24'b010010100000000001001110;
			 rom[567] = 24'b010101010111001100000000;
			 rom[568] = 24'b010010100000000001001110;
			 rom[569] = 24'b001010101011100110000000;
			 rom[570] = 24'b000000000000000000000000;
			 rom[571] = 24'b110101010100011010000000;
			 rom[572] = 24'b101101011111111110110010;
			 rom[573] = 24'b101010101000110100000000;
			 rom[574] = 24'b101101011111111110110010;
			 rom[575] = 24'b110101010100011010000000;
			 rom[576] = 24'b000000000000000000000000;
			 rom[577] = 24'b001010101011100110000000;
			 rom[578] = 24'b010010100000000001001110;
			 rom[579] = 24'b010101010111001100000000;
			 rom[580] = 24'b010010100000000001001110;
			 rom[581] = 24'b001010101011100110000000;
			 rom[582] = 24'b000000000000000000000000;
			 rom[583] = 24'b110101010100011010000000;
			 rom[584] = 24'b101101011111111110110010;
			 rom[585] = 24'b101010101000110100000000;
			 rom[586] = 24'b101101011111111110110010;
			 rom[587] = 24'b110101010100011010000000;
			 rom[588] = 24'b000000000000000000000000;
			 rom[589] = 24'b001010101011100110000000;
			 rom[590] = 24'b010010100000000001001110;
			 rom[591] = 24'b010101010111001100000000;
			 rom[592] = 24'b010010100000000001001110;
			 rom[593] = 24'b001010101011100110000000;
			 rom[594] = 24'b000000000000000000000000;
			 rom[595] = 24'b110101010100011010000000;
			 rom[596] = 24'b101101011111111110110010;
			 rom[597] = 24'b101010101000110100000000;
			 rom[598] = 24'b101101011111111110110010;
			 rom[599] = 24'b110101010100011010000000;
			 rom[600] = 24'b000000000000000000000000;
			 rom[601] = 24'b001010101011100110000000;
			 rom[602] = 24'b010010100000000001001110;
			 rom[603] = 24'b010101010111001100000000;
			 rom[604] = 24'b010010100000000001001110;
			 rom[605] = 24'b001010101011100110000000;
			 rom[606] = 24'b000000000000000000000000;
			 rom[607] = 24'b110101010100011010000000;
			 rom[608] = 24'b101101011111111110110010;
			 rom[609] = 24'b101010101000110100000000;
			 rom[610] = 24'b101101011111111110110010;
			 rom[611] = 24'b110101010100011010000000;
			 rom[612] = 24'b000000000000000000000000;
			 rom[613] = 24'b001010101011100110000000;
			 rom[614] = 24'b010010100000000001001110;
			 rom[615] = 24'b010101010111001100000000;
			 rom[616] = 24'b010010100000000001001110;
			 rom[617] = 24'b001010101011100110000000;
			 rom[618] = 24'b000000000000000000000000;
			 rom[619] = 24'b110101010100011010000000;
			 rom[620] = 24'b101101011111111110110010;
			 rom[621] = 24'b101010101000110100000000;
			 rom[622] = 24'b101101011111111110110010;
			 rom[623] = 24'b110101010100011010000000;
			 rom[624] = 24'b000000000000000000000000;
			 rom[625] = 24'b001010101011100110000000;
			 rom[626] = 24'b010010100000000001001110;
			 rom[627] = 24'b010101010111001100000000;
			 rom[628] = 24'b010010100000000001001110;
			 rom[629] = 24'b001010101011100110000000;
			 rom[630] = 24'b000000000000000000000000;
			 rom[631] = 24'b110101010100011010000000;
			 rom[632] = 24'b101101011111111110110010;
			 rom[633] = 24'b101010101000110100000000;
			 rom[634] = 24'b101101011111111110110010;
			 rom[635] = 24'b110101010100011010000000;
			 rom[636] = 24'b000000000000000000000000;
			 rom[637] = 24'b001010101011100110000000;
			 rom[638] = 24'b010010100000000001001110;
			 rom[639] = 24'b010101010111001100000000;
			 rom[640] = 24'b010010100000000001001110;
			 rom[641] = 24'b001010101011100110000000;
			 rom[642] = 24'b000000000000000000000000;
			 rom[643] = 24'b110101010100011010000000;
			 rom[644] = 24'b101101011111111110110010;
			 rom[645] = 24'b101010101000110100000000;
			 rom[646] = 24'b101101011111111110110010;
			 rom[647] = 24'b110101010100011010000000;
			 rom[648] = 24'b000000000000000000000000;
			 rom[649] = 24'b001010101011100110000000;
			 rom[650] = 24'b010010100000000001001110;
			 rom[651] = 24'b010101010111001100000000;
			 rom[652] = 24'b010010100000000001001110;
			 rom[653] = 24'b001010101011100110000000;
			 rom[654] = 24'b000000000000000000000000;
			 rom[655] = 24'b110101010100011010000000;
			 rom[656] = 24'b101101011111111110110010;
			 rom[657] = 24'b101010101000110100000000;
			 rom[658] = 24'b101101011111111110110010;
			 rom[659] = 24'b110101010100011010000000;
			 rom[660] = 24'b000000000000000000000000;
			 rom[661] = 24'b001010101011100110000000;
			 rom[662] = 24'b010010100000000001001110;
			 rom[663] = 24'b010101010111001100000000;
			 rom[664] = 24'b010010100000000001001110;
			 rom[665] = 24'b001010101011100110000000;
			 rom[666] = 24'b000000000000000000000000;
			 rom[667] = 24'b110101010100011010000000;
			 rom[668] = 24'b101101011111111110110010;
			 rom[669] = 24'b101010101000110100000000;
			 rom[670] = 24'b101101011111111110110010;
			 rom[671] = 24'b110101010100011010000000;
			 rom[672] = 24'b000000000000000000000000;
			 rom[673] = 24'b001010101011100110000000;
			 rom[674] = 24'b010010100000000001001110;
			 rom[675] = 24'b010101010111001100000000;
			 rom[676] = 24'b010010100000000001001110;
			 rom[677] = 24'b001010101011100110000000;
			 rom[678] = 24'b000000000000000000000000;
			 rom[679] = 24'b110101010100011010000000;
			 rom[680] = 24'b101101011111111110110010;
			 rom[681] = 24'b101010101000110100000000;
			 rom[682] = 24'b101101011111111110110010;
			 rom[683] = 24'b110101010100011010000000;
			 rom[684] = 24'b000000000000000000000000;
			 rom[685] = 24'b001010101011100110000000;
			 rom[686] = 24'b010010100000000001001110;
			 rom[687] = 24'b010101010111001100000000;
			 rom[688] = 24'b010010100000000001001110;
			 rom[689] = 24'b001010101011100110000000;
			 rom[690] = 24'b000000000000000000000000;
			 rom[691] = 24'b110101010100011010000000;
			 rom[692] = 24'b101101011111111110110010;
			 rom[693] = 24'b101010101000110100000000;
			 rom[694] = 24'b101101011111111110110010;
			 rom[695] = 24'b110101010100011010000000;
			 rom[696] = 24'b000000000000000000000000;
			 rom[697] = 24'b001010101011100110000000;
			 rom[698] = 24'b010010100000000001001110;
			 rom[699] = 24'b010101010111001100000000;
			 rom[700] = 24'b010010100000000001001110;
			 rom[701] = 24'b001010101011100110000000;
			 rom[702] = 24'b000000000000000000000000;
			 rom[703] = 24'b110101010100011010000000;
			 rom[704] = 24'b101101011111111110110010;
			 rom[705] = 24'b101010101000110100000000;
			 rom[706] = 24'b101101011111111110110010;
			 rom[707] = 24'b110101010100011010000000;
			 rom[708] = 24'b000000000000000000000000;
			 rom[709] = 24'b001010101011100110000000;
			 rom[710] = 24'b010010100000000001001110;
			 rom[711] = 24'b010101010111001100000000;
			 rom[712] = 24'b010010100000000001001110;
			 rom[713] = 24'b001010101011100110000000;
			 rom[714] = 24'b000000000000000000000000;
			 rom[715] = 24'b110101010100011010000000;
			 rom[716] = 24'b101101011111111110110010;
			 rom[717] = 24'b101010101000110100000000;
			 rom[718] = 24'b101101011111111110110010;
			 rom[719] = 24'b110101010100011010000000;
			 rom[720] = 24'b000000000000000000000000;
			 rom[721] = 24'b001010101011100110000000;
			 rom[722] = 24'b010010100000000001001110;
			 rom[723] = 24'b010101010111001100000000;
			 rom[724] = 24'b010010100000000001001110;
			 rom[725] = 24'b001010101011100110000000;
			 rom[726] = 24'b000000000000000000000000;
			 rom[727] = 24'b110101010100011010000000;
			 rom[728] = 24'b101101011111111110110010;
			 rom[729] = 24'b101010101000110100000000;
			 rom[730] = 24'b101101011111111110110010;
			 rom[731] = 24'b110101010100011010000000;
			 rom[732] = 24'b000000000000000000000000;
			 rom[733] = 24'b001010101011100110000000;
			 rom[734] = 24'b010010100000000001001110;
			 rom[735] = 24'b010101010111001100000000;
			 rom[736] = 24'b010010100000000001001110;
			 rom[737] = 24'b001010101011100110000000;
			 rom[738] = 24'b000000000000000000000000;
			 rom[739] = 24'b110101010100011010000000;
			 rom[740] = 24'b101101011111111110110010;
			 rom[741] = 24'b101010101000110100000000;
			 rom[742] = 24'b101101011111111110110010;
			 rom[743] = 24'b110101010100011010000000;
			 rom[744] = 24'b000000000000000000000000;
			 rom[745] = 24'b001010101011100110000000;
			 rom[746] = 24'b010010100000000001001110;
			 rom[747] = 24'b010101010111001100000000;
			 rom[748] = 24'b010010100000000001001110;
			 rom[749] = 24'b001010101011100110000000;
			 rom[750] = 24'b000000000000000000000000;
			 rom[751] = 24'b110101010100011010000000;
			 rom[752] = 24'b101101011111111110110010;
			 rom[753] = 24'b101010101000110100000000;
			 rom[754] = 24'b101101011111111110110010;
			 rom[755] = 24'b110101010100011010000000;
			 rom[756] = 24'b000000000000000000000000;
			 rom[757] = 24'b001010101011100110000000;
			 rom[758] = 24'b010010100000000001001110;
			 rom[759] = 24'b010101010111001100000000;
			 rom[760] = 24'b010010100000000001001110;
			 rom[761] = 24'b001010101011100110000000;
			 rom[762] = 24'b000000000000000000000000;
			 rom[763] = 24'b110101010100011010000000;
			 rom[764] = 24'b101101011111111110110010;
			 rom[765] = 24'b101010101000110100000000;
			 rom[766] = 24'b101101011111111110110010;
			 rom[767] = 24'b110101010100011010000000;
			 rom[768] = 24'b000000000000000000000000;
			 rom[769] = 24'b001010101011100110000000;
			 rom[770] = 24'b010010100000000001001110;
			 rom[771] = 24'b010101010111001100000000;
			 rom[772] = 24'b010010100000000001001110;
			 rom[773] = 24'b001010101011100110000000;
			 rom[774] = 24'b000000000000000000000000;
			 rom[775] = 24'b110101010100011010000000;
			 rom[776] = 24'b101101011111111110110010;
			 rom[777] = 24'b101010101000110100000000;
			 rom[778] = 24'b101101011111111110110010;
			 rom[779] = 24'b110101010100011010000000;
			 rom[780] = 24'b000000000000000000000000;
			 rom[781] = 24'b001010101011100110000000;
			 rom[782] = 24'b010010100000000001001110;
			 rom[783] = 24'b010101010111001100000000;
			 rom[784] = 24'b010010100000000001001110;
			 rom[785] = 24'b001010101011100110000000;
			 rom[786] = 24'b000000000000000000000000;
			 rom[787] = 24'b110101010100011010000000;
			 rom[788] = 24'b101101011111111110110010;
			 rom[789] = 24'b101010101000110100000000;
			 rom[790] = 24'b101101011111111110110010;
			 rom[791] = 24'b110101010100011010000000;
			 rom[792] = 24'b000000000000000000000000;
			 rom[793] = 24'b001010101011100110000000;
			 rom[794] = 24'b010010100000000001001110;
			 rom[795] = 24'b010101010111001100000000;
			 rom[796] = 24'b010010100000000001001110;
			 rom[797] = 24'b001010101011100110000000;
			 rom[798] = 24'b000000000000000000000000;
			 rom[799] = 24'b110101010100011010000000;
			 rom[800] = 24'b101101011111111110110010;
			 rom[801] = 24'b101010101000110100000000;
			 rom[802] = 24'b101101011111111110110010;
			 rom[803] = 24'b110101010100011010000000;
			 rom[804] = 24'b000000000000000000000000;
			 rom[805] = 24'b001010101011100110000000;
			 rom[806] = 24'b010010100000000001001110;
			 rom[807] = 24'b010101010111001100000000;
			 rom[808] = 24'b010010100000000001001110;
			 rom[809] = 24'b001010101011100110000000;
			 rom[810] = 24'b000000000000000000000000;
			 rom[811] = 24'b110101010100011010000000;
			 rom[812] = 24'b101101011111111110110010;
			 rom[813] = 24'b101010101000110100000000;
			 rom[814] = 24'b101101011111111110110010;
			 rom[815] = 24'b110101010100011010000000;
			 rom[816] = 24'b000000000000000000000000;
			 rom[817] = 24'b001010101011100110000000;
			 rom[818] = 24'b010010100000000001001110;
			 rom[819] = 24'b010101010111001100000000;
			 rom[820] = 24'b010010100000000001001110;
			 rom[821] = 24'b001010101011100110000000;
			 rom[822] = 24'b000000000000000000000000;
			 rom[823] = 24'b110101010100011010000000;
			 rom[824] = 24'b101101011111111110110010;
			 rom[825] = 24'b101010101000110100000000;
			 rom[826] = 24'b101101011111111110110010;
			 rom[827] = 24'b110101010100011010000000;
			 rom[828] = 24'b000000000000000000000000;
			 rom[829] = 24'b001010101011100110000000;
			 rom[830] = 24'b010010100000000001001110;
			 rom[831] = 24'b010101010111001100000000;
			 rom[832] = 24'b010010100000000001001110;
			 rom[833] = 24'b001010101011100110000000;
			 rom[834] = 24'b000000000000000000000000;
			 rom[835] = 24'b110101010100011010000000;
			 rom[836] = 24'b101101011111111110110010;
			 rom[837] = 24'b101010101000110100000000;
			 rom[838] = 24'b101101011111111110110010;
			 rom[839] = 24'b110101010100011010000000;
			 rom[840] = 24'b000000000000000000000000;
			 rom[841] = 24'b001010101011100110000000;
			 rom[842] = 24'b010010100000000001001110;
			 rom[843] = 24'b010101010111001100000000;
			 rom[844] = 24'b010010100000000001001110;
			 rom[845] = 24'b001010101011100110000000;
			 rom[846] = 24'b000000000000000000000000;
			 rom[847] = 24'b110101010100011010000000;
			 rom[848] = 24'b101101011111111110110010;
			 rom[849] = 24'b101010101000110100000000;
			 rom[850] = 24'b101101011111111110110010;
			 rom[851] = 24'b110101010100011010000000;
			 rom[852] = 24'b000000000000000000000000;
			 rom[853] = 24'b001010101011100110000000;
			 rom[854] = 24'b010010100000000001001110;
			 rom[855] = 24'b010101010111001100000000;
			 rom[856] = 24'b010010100000000001001110;
			 rom[857] = 24'b001010101011100110000000;
			 rom[858] = 24'b000000000000000000000000;
			 rom[859] = 24'b110101010100011010000000;
			 rom[860] = 24'b101101011111111110110010;
			 rom[861] = 24'b101010101000110100000000;
			 rom[862] = 24'b101101011111111110110010;
			 rom[863] = 24'b110101010100011010000000;
			 rom[864] = 24'b000000000000000000000000;
			 rom[865] = 24'b001010101011100110000000;
			 rom[866] = 24'b010010100000000001001110;
			 rom[867] = 24'b010101010111001100000000;
			 rom[868] = 24'b010010100000000001001110;
			 rom[869] = 24'b001010101011100110000000;
			 rom[870] = 24'b000000000000000000000000;
			 rom[871] = 24'b110101010100011010000000;
			 rom[872] = 24'b101101011111111110110010;
			 rom[873] = 24'b101010101000110100000000;
			 rom[874] = 24'b101101011111111110110010;
			 rom[875] = 24'b110101010100011010000000;
			 rom[876] = 24'b000000000000000000000000;
			 rom[877] = 24'b001010101011100110000000;
			 rom[878] = 24'b010010100000000001001110;
			 rom[879] = 24'b010101010111001100000000;
			 rom[880] = 24'b010010100000000001001110;
			 rom[881] = 24'b001010101011100110000000;
			 rom[882] = 24'b000000000000000000000000;
			 rom[883] = 24'b110101010100011010000000;
			 rom[884] = 24'b101101011111111110110010;
			 rom[885] = 24'b101010101000110100000000;
			 rom[886] = 24'b101101011111111110110010;
			 rom[887] = 24'b110101010100011010000000;
			 rom[888] = 24'b000000000000000000000000;
			 rom[889] = 24'b001010101011100110000000;
			 rom[890] = 24'b010010100000000001001110;
			 rom[891] = 24'b010101010111001100000000;
			 rom[892] = 24'b010010100000000001001110;
			 rom[893] = 24'b001010101011100110000000;
			 rom[894] = 24'b000000000000000000000000;
			 rom[895] = 24'b110101010100011010000000;
			 rom[896] = 24'b101101011111111110110010;
			 rom[897] = 24'b101010101000110100000000;
			 rom[898] = 24'b101101011111111110110010;
			 rom[899] = 24'b110101010100011010000000;
			 rom[900] = 24'b000000000000000000000000;
			 rom[901] = 24'b001010101011100110000000;
			 rom[902] = 24'b010010100000000001001110;
			 rom[903] = 24'b010101010111001100000000;
			 rom[904] = 24'b010010100000000001001110;
			 rom[905] = 24'b001010101011100110000000;
			 rom[906] = 24'b000000000000000000000000;
			 rom[907] = 24'b110101010100011010000000;
			 rom[908] = 24'b101101011111111110110010;
			 rom[909] = 24'b101010101000110100000000;
			 rom[910] = 24'b101101011111111110110010;
			 rom[911] = 24'b110101010100011010000000;
			 rom[912] = 24'b000000000000000000000000;
			 rom[913] = 24'b001010101011100110000000;
			 rom[914] = 24'b010010100000000001001110;
			 rom[915] = 24'b010101010111001100000000;
			 rom[916] = 24'b010010100000000001001110;
			 rom[917] = 24'b001010101011100110000000;
			 rom[918] = 24'b000000000000000000000000;
			 rom[919] = 24'b110101010100011010000000;
			 rom[920] = 24'b101101011111111110110010;
			 rom[921] = 24'b101010101000110100000000;
			 rom[922] = 24'b101101011111111110110010;
			 rom[923] = 24'b110101010100011010000000;
			 rom[924] = 24'b000000000000000000000000;
			 rom[925] = 24'b001010101011100110000000;
			 rom[926] = 24'b010010100000000001001110;
			 rom[927] = 24'b010101010111001100000000;
			 rom[928] = 24'b010010100000000001001110;
			 rom[929] = 24'b001010101011100110000000;
			 rom[930] = 24'b000000000000000000000000;
			 rom[931] = 24'b110101010100011010000000;
			 rom[932] = 24'b101101011111111110110010;
			 rom[933] = 24'b101010101000110100000000;
			 rom[934] = 24'b101101011111111110110010;
			 rom[935] = 24'b110101010100011010000000;
			 rom[936] = 24'b000000000000000000000000;
			 rom[937] = 24'b001010101011100110000000;
			 rom[938] = 24'b010010100000000001001110;
			 rom[939] = 24'b010101010111001100000000;
			 rom[940] = 24'b010010100000000001001110;
			 rom[941] = 24'b001010101011100110000000;
			 rom[942] = 24'b000000000000000000000000;
			 rom[943] = 24'b110101010100011010000000;
			 rom[944] = 24'b101101011111111110110010;
			 rom[945] = 24'b101010101000110100000000;
			 rom[946] = 24'b101101011111111110110010;
			 rom[947] = 24'b110101010100011010000000;
			 rom[948] = 24'b000000000000000000000000;
			 rom[949] = 24'b001010101011100110000000;
			 rom[950] = 24'b010010100000000001001110;
			 rom[951] = 24'b010101010111001100000000;
			 rom[952] = 24'b010010100000000001001110;
			 rom[953] = 24'b001010101011100110000000;
			 rom[954] = 24'b000000000000000000000000;
			 rom[955] = 24'b110101010100011010000000;
			 rom[956] = 24'b101101011111111110110010;
			 rom[957] = 24'b101010101000110100000000;
			 rom[958] = 24'b101101011111111110110010;
			 rom[959] = 24'b110101010100011010000000;
		 end 

	 always @(posedge(clk))
		 begin 
			 if(reset) 
				 begin 
					 data_out <= 24'b0; 
					 i <= 16'b0; 
					 counter <= 16'b0; 
				 end 
			 else 
				 begin 
					 if(counter == 16'd2083) 
						 begin 
							 data_out <= rom[i]; 
							 counter <=16'b0; 
							 if(i == 959) i <= 0; 
							 else i <= i + 1; 
						 end 
					 else counter <= counter + 16'd1; 
				 end 
		 end 

endmodule
