//////////////////////////////////////////////////////////////////////////////////
// Kolo Naukowe Systemow Scalonych
// 10.2017
// 
// Modul: gen_sinus
// Projekt: Adaptacyjne filtry cyfrowe do kondycjonowania sygnalow biomedycznych 
// Model urzadzenia: Nexys Video Artix 7 (XC7A200T-1SBG484C)
// 
// Wersja: 0.1
//////////////////////////////////////////////////////////////////////////////////


module gen_sinus(
    output reg signed [23:0] data_out,
    input clk,
    input reset
    );
    
    reg signed [23:0] rom [0:39];
    reg [8:0] i;
    reg [15:0] counter;//50000 * 40pr�bek = 2 000 000 ; zegar 100mhz => 50hz

    always @(reset)
        begin
        rom[0] = 24'b000000000000000000000000;
        rom[1] = 24'b000011010101111000000001;
        rom[2] = 24'b000110100110011110111111;
        rom[3] = 24'b001001101100101100001011;
        rom[4] = 24'b001100100011100111001101;
        rom[5] = 24'b001111000110101111110110;
        rom[6] = 24'b010001010010000100111111;
        rom[7] = 24'b010011000010001011000101;
        rom[8] = 24'b010100010100010001011100;
        rom[9] = 24'b010101000110010110101111;
        rom[10] = 24'b010101010111001100000000;
        rom[11] = 24'b010101000110010110101111;
        rom[12] = 24'b010100010100010001011100;
        rom[13] = 24'b010011000010001011000101;
        rom[14] = 24'b010001010010000100111111;
        rom[15] = 24'b001111000110101111110110;
        rom[16] = 24'b001100100011100111001101;
        rom[17] = 24'b001001101100101100001011;
        rom[18] = 24'b000110100110011110111111;
        rom[19] = 24'b000011010101111000000001;
        rom[20] = 24'b000000000000000000000000;
        rom[21] = 24'b111100101010000111111111;
        rom[22] = 24'b111001011001100001000001;
        rom[23] = 24'b110110010011010011110101;
        rom[24] = 24'b110011011100011000110011;
        rom[25] = 24'b110000111001010000001010;
        rom[26] = 24'b101110101101111011000001;
        rom[27] = 24'b101100111101110100111011;
        rom[28] = 24'b101011101011101110100100;
        rom[29] = 24'b101010111001101001010001;
        rom[30] = 24'b101010101000110100000000;
        rom[31] = 24'b101010111001101001010001;
        rom[32] = 24'b101011101011101110100100;
        rom[33] = 24'b101100111101110100111011;
        rom[34] = 24'b101110101101111011000001;
        rom[35] = 24'b110000111001010000001010;
        rom[36] = 24'b110011011100011000110011;
        rom[37] = 24'b110110010011010011110101;
        rom[38] = 24'b111001011001100001000001;
        rom[39] = 24'b111100101010000111111111;

        end
        
        always @(posedge(clk))
            begin
                if(reset)
                    begin
                        data_out <= 24'b0;
                        i <= 9'b0;
                        counter <= 16'b0;
                    end
                else
                    begin
                        if(counter == 16'd50000)
                            begin
                                data_out <= rom[i];
                                counter <= 16'b0;
                                if(i == 39) i <= 0;
                                else i <= i + 1;
                            end
                        else counter <= counter + 16'd1;
                    end
            end
            
endmodule
