//////////////////////////////////////////////////////////////////////////////////
// Kolo Naukowe Systemow Scalonych
// 10.2017
// 
// Modul: gen_ekg_zabrudzony
// Projekt: Adaptacyjne filtry cyfrowe do kondycjonowania sygnalow biomedycznych 
// Model urzadzenia: Nexys Video Artix 7 (XC7A200T-1SBG484C)
// 
// Wersja: 0.1
//////////////////////////////////////////////////////////////////////////////////


module gen_ekg_zabrudzony(
    output reg signed [23:0] data_out,
    input clk,
    input reset
    );
    
    reg signed [23:0] rom [0:3599];
    reg [15:0] i;
    reg [19:0] counter;//360000 * 3600pr�bek /13 okresow= 100 000 000 ; zegar 100mhz => 1hz

    always @(reset)
        begin
        rom[0] = 24'b000100000000010110010000;
        rom[1] = 24'b000100110111101010100000;
        rom[2] = 24'b000100101111000110100111;
        rom[3] = 24'b000011110000100011001111;
        rom[4] = 24'b000011000100001111010110;
        rom[5] = 24'b000011011101010101101101;
        rom[6] = 24'b000100011110110111011000;
        rom[7] = 24'b000100111101001001101000;
        rom[8] = 24'b000100100001011011100001;
        rom[9] = 24'b000011011010000100100111;
        rom[10] = 24'b000011000110111111100100;
        rom[11] = 24'b000011111000100101100011;
        rom[12] = 24'b000100101101111000011010;
        rom[13] = 24'b000100101101011101100100;
        rom[14] = 24'b000011101110011011001011;
        rom[15] = 24'b000010110110101111100110;
        rom[16] = 24'b000011001000000001100111;
        rom[17] = 24'b000100000110100111000110;
        rom[18] = 24'b000100110001001011010000;
        rom[19] = 24'b000100010101010000100110;
        rom[20] = 24'b000011001010011101110111;
        rom[21] = 24'b000010110100010011010110;
        rom[22] = 24'b000011011111110001101011;
        rom[23] = 24'b000100100001010000010100;
        rom[24] = 24'b000100110000010100101010;
        rom[25] = 24'b000011111111111010010011;
        rom[26] = 24'b000011000010000111000100;
        rom[27] = 24'b000010111111001101110111;
        rom[28] = 24'b000011110111111011010001;
        rom[29] = 24'b000100010001001101001000;
        rom[30] = 24'b000011110111110011010111;
        rom[31] = 24'b000010101100100000101101;
        rom[32] = 24'b000010010000111110000110;
        rom[33] = 24'b000010111000011001011111;
        rom[34] = 24'b000011101111101000000111;
        rom[35] = 24'b000011111000001100000000;
        rom[36] = 24'b000011000000110111101111;
        rom[37] = 24'b000010001110011011111111;
        rom[38] = 24'b000010011011111000011000;
        rom[39] = 24'b000011010101100011010000;
        rom[40] = 24'b000011111100111110101001;
        rom[41] = 24'b000011011100100011100010;
        rom[42] = 24'b000010011011000001111000;
        rom[43] = 24'b000001111100101111100111;
        rom[44] = 24'b000010100100101010111110;
        rom[45] = 24'b000011100111001001011000;
        rom[46] = 24'b000011110000011101011011;
        rom[47] = 24'b000010110111100010101100;
        rom[48] = 24'b000010000111001000010101;
        rom[49] = 24'b000010001110110111111011;
        rom[50] = 24'b000011001011011110000100;
        rom[51] = 24'b000011111001011000101001;
        rom[52] = 24'b000011100011001110001000;
        rom[53] = 24'b000010011000011011011001;
        rom[54] = 24'b000001111100100000110000;
        rom[55] = 24'b000010011010110111101001;
        rom[56] = 24'b000011100101101010011000;
        rom[57] = 24'b000011110100100000001001;
        rom[58] = 24'b000010111111010000110100;
        rom[59] = 24'b000001111011010101111011;
        rom[60] = 24'b000001110110000010100101;
        rom[61] = 24'b000010101000111001001100;
        rom[62] = 24'b000011010000101110001011;
        rom[63] = 24'b000010110110010100011000;
        rom[64] = 24'b000001110110010010001110;
        rom[65] = 24'b000001000100100101110111;
        rom[66] = 24'b000001001010011101101000;
        rom[67] = 24'b000001111101010101110010;
        rom[68] = 24'b000010010110011100001001;
        rom[69] = 24'b000010000111011011010000;
        rom[70] = 24'b000001110111010000101000;
        rom[71] = 24'b000010100100011010001111;
        rom[72] = 24'b000100100100111110000000;
        rom[73] = 24'b000110111001000011110000;
        rom[74] = 24'b001000101101000000100111;
        rom[75] = 24'b001001100110000101011111;
        rom[76] = 24'b001010000111111001100110;
        rom[77] = 24'b001010111110010010111101;
        rom[78] = 24'b001011011011001100111000;
        rom[79] = 24'b001010000001110110111000;
        rom[80] = 24'b000110101111000010000001;
        rom[81] = 24'b000011001011011011000111;
        rom[82] = 24'b000001011011100100100100;
        rom[83] = 24'b000001101101011011010011;
        rom[84] = 24'b000010101100011111001010;
        rom[85] = 24'b000011000100011110110100;
        rom[86] = 24'b000010011011011010101011;
        rom[87] = 24'b000001101101100000000110;
        rom[88] = 24'b000001111100010101110111;
        rom[89] = 24'b000010111000011111000110;
        rom[90] = 24'b000011100011000011010000;
        rom[91] = 24'b000011000010010000000110;
        rom[92] = 24'b000010000110000110110111;
        rom[93] = 24'b000001110100110100110110;
        rom[94] = 24'b000010100000010011001011;
        rom[95] = 24'b000011010101100100100100;
        rom[96] = 24'b000011010101111111011010;
        rom[97] = 24'b000010100011001000110011;
        rom[98] = 24'b000001100101010101100100;
        rom[99] = 24'b000001111000011010100111;
        rom[100] = 24'b000010111010111001000001;
        rom[101] = 24'b000011100000011000001000;
        rom[102] = 24'b000011000100100010000111;
        rom[103] = 24'b000010000101011100101101;
        rom[104] = 24'b000001101001111010000110;
        rom[105] = 24'b000010010110001101111111;
        rom[106] = 24'b000011001101011100100111;
        rom[107] = 24'b000011010001001000000000;
        rom[108] = 24'b000010100011100100101111;
        rom[109] = 24'b000001110001001000111111;
        rom[110] = 24'b000010000011011101111000;
        rom[111] = 24'b000010111010101100100000;
        rom[112] = 24'b000011100111000000011001;
        rom[113] = 24'b000011001001000001100010;
        rom[114] = 24'b000010000010100111010111;
        rom[115] = 24'b000001100110110001010111;
        rom[116] = 24'b000010001100010000011110;
        rom[117] = 24'b000011001001110110011000;
        rom[118] = 24'b000011010011001010011011;
        rom[119] = 24'b000010011111001000001100;
        rom[120] = 24'b000001101100010001100101;
        rom[121] = 24'b000001110100000001001011;
        rom[122] = 24'b000010110000100111010100;
        rom[123] = 24'b000011100000111110001001;
        rom[124] = 24'b000011001000010111011000;
        rom[125] = 24'b000010000010011101001001;
        rom[126] = 24'b000001101011011011000000;
        rom[127] = 24'b000010001110101010011001;
        rom[128] = 24'b000011001101001111111000;
        rom[129] = 24'b000011100000111110001001;
        rom[130] = 24'b000010101110001011000100;
        rom[131] = 24'b000001110001100100111011;
        rom[132] = 24'b000001101100010001100101;
        rom[133] = 24'b000010101011010101011100;
        rom[134] = 24'b000011011010011111001011;
        rom[135] = 24'b000011000111011010001000;
        rom[136] = 24'b000010000100111011101110;
        rom[137] = 24'b000001011111011100100111;
        rom[138] = 24'b000010000000001011001000;
        rom[139] = 24'b000011001001000001100010;
        rom[140] = 24'b000011100111000000011001;
        rom[141] = 24'b000010110011010111110000;
        rom[142] = 24'b000001110111010000101000;
        rom[143] = 24'b000001100111010111111111;
        rom[144] = 24'b000010100110000001000000;
        rom[145] = 24'b000011011010111001000000;
        rom[146] = 24'b000011010010010101000111;
        rom[147] = 24'b000010001110111001001111;
        rom[148] = 24'b000001100010100101010110;
        rom[149] = 24'b000001110110110011001101;
        rom[150] = 24'b000010111111101001101000;
        rom[151] = 24'b000011011101111011111000;
        rom[152] = 24'b000010111000011100110001;
        rom[153] = 24'b000001111010110110110111;
        rom[154] = 24'b000001100010111001010100;
        rom[155] = 24'b000010010110111011100011;
        rom[156] = 24'b000011010011100011001010;
        rom[157] = 24'b000011010101100100100100;
        rom[158] = 24'b000010011000111110011011;
        rom[159] = 24'b000001101000100111100110;
        rom[160] = 24'b000001110101000001000111;
        rom[161] = 24'b000010110011100110100110;
        rom[162] = 24'b000011010110110110000000;
        rom[163] = 24'b000010111000011111000110;
        rom[164] = 24'b000001110111011101010111;
        rom[165] = 24'b000001101000100111100110;
        rom[166] = 24'b000010010001101001101011;
        rom[167] = 24'b000011001001010111010100;
        rom[168] = 24'b000011001100001110011010;
        rom[169] = 24'b000010010010000011000011;
        rom[170] = 24'b000001011011100100100100;
        rom[171] = 24'b000001101100001101010111;
        rom[172] = 24'b000010100111010111000001;
        rom[173] = 24'b000011000111111101101000;
        rom[174] = 24'b000010110001000000000111;
        rom[175] = 24'b000001110100010110111101;
        rom[176] = 24'b000001011101101100110110;
        rom[177] = 24'b000010000111100100011111;
        rom[178] = 24'b000010111110110011000111;
        rom[179] = 24'b000011000111010111000000;
        rom[180] = 24'b000010010100111011001111;
        rom[181] = 24'b000001011101100110111111;
        rom[182] = 24'b000001101000100111001000;
        rom[183] = 24'b000010100111001010100000;
        rom[184] = 24'b000011010001000010001001;
        rom[185] = 24'b000010110101011111100010;
        rom[186] = 24'b000001111011010010100111;
        rom[187] = 24'b000001101001001101100111;
        rom[188] = 24'b000010010011100101001110;
        rom[189] = 24'b000011010011100111011000;
        rom[190] = 24'b000011011100111011011011;
        rom[191] = 24'b000010100110011100111100;
        rom[192] = 24'b000001111000011110110101;
        rom[193] = 24'b000010000010101010101011;
        rom[194] = 24'b000010111111010000110100;
        rom[195] = 24'b000011110100100000001001;
        rom[196] = 24'b000011011110010101101000;
        rom[197] = 24'b000010011111110000001001;
        rom[198] = 24'b000001111110111101000000;
        rom[199] = 24'b000010100111000100111001;
        rom[200] = 24'b000011110001110111101000;
        rom[201] = 24'b000100001000000010001001;
        rom[202] = 24'b000011010111101011010100;
        rom[203] = 24'b000010010011110000011011;
        rom[204] = 24'b000010010101110001110101;
        rom[205] = 24'b000011010100110101101100;
        rom[206] = 24'b000100010000001100101011;
        rom[207] = 24'b000011111010101011011000;
        rom[208] = 24'b000010111010101001001110;
        rom[209] = 24'b000010001101110101010111;
        rom[210] = 24'b000010101100000111101000;
        rom[211] = 24'b000011110100111110000010;
        rom[212] = 24'b000100001001001011111001;
        rom[213] = 24'b000011011010011011110000;
        rom[214] = 24'b000010100000110000111000;
        rom[215] = 24'b000010010011010100011111;
        rom[216] = 24'b000011001101000101000000;
        rom[217] = 24'b000100000100011001010000;
        rom[218] = 24'b000011110100100000100111;
        rom[219] = 24'b000010111000011001011111;
        rom[220] = 24'b000010001100000101100110;
        rom[221] = 24'b000010100010101111101101;
        rom[222] = 24'b000011100001110101001000;
        rom[223] = 24'b000100000010100011101000;
        rom[224] = 24'b000011011101000100100001;
        rom[225] = 24'b000010010101101101100111;
        rom[226] = 24'b000010000101000100110100;
        rom[227] = 24'b000010110100001110100011;
        rom[228] = 24'b000011110101101110101010;
        rom[229] = 24'b000011110101010011110100;
        rom[230] = 24'b000010111101100110001011;
        rom[231] = 24'b000010000011011110010110;
        rom[232] = 24'b000010010111001100100111;
        rom[233] = 24'b000011010101110010000110;
        rom[234] = 24'b000011111101111010000000;
        rom[235] = 24'b000011011010101010100110;
        rom[236] = 24'b000010011110100001010111;
        rom[237] = 24'b000010001000010110110110;
        rom[238] = 24'b000010110001011000111011;
        rom[239] = 24'b000011101011100010110100;
        rom[240] = 24'b000011110011010010011010;
        rom[241] = 24'b000010111011100011010011;
        rom[242] = 24'b000010000010101000100100;
        rom[243] = 24'b000010010011010001010111;
        rom[244] = 24'b000011001001100010100001;
        rom[245] = 24'b000011110001011101111000;
        rom[246] = 24'b000011010000101111011000;
        rom[247] = 24'b000010010100000110001101;
        rom[248] = 24'b000001111000100011100110;
        rom[249] = 24'b000010011111111110111111;
        rom[250] = 24'b000011011110100010010111;
        rom[251] = 24'b000011101001100010100000;
        rom[252] = 24'b000010110111000110110000;
        rom[253] = 24'b000010000100101010111111;
        rom[254] = 24'b000010001101001110111000;
        rom[255] = 24'b000011001001010110000000;
        rom[256] = 24'b000011110011001101101001;
        rom[257] = 24'b000011010010110010100010;
        rom[258] = 24'b000010011011000001111000;
        rom[259] = 24'b000001111010010011010111;
        rom[260] = 24'b000010011111110010011110;
        rom[261] = 24'b000011011101011000011000;
        rom[262] = 24'b000011101001001000101011;
        rom[263] = 24'b000010101101110001101100;
        rom[264] = 24'b000001111010111011000101;
        rom[265] = 24'b000010000010101010101011;
        rom[266] = 24'b000011000100001001010100;
        rom[267] = 24'b000011101010101111001001;
        rom[268] = 24'b000011001111101100001000;
        rom[269] = 24'b000010001100001110001001;
        rom[270] = 24'b000001110000010011100000;
        rom[271] = 24'b000010011010110111101001;
        rom[272] = 24'b000011011001011101001000;
        rom[273] = 24'b000011101010101111001001;
        rom[274] = 24'b000010110101011111110100;
        rom[275] = 24'b000001110100000001001011;
        rom[276] = 24'b000001110011100110010101;
        rom[277] = 24'b000010110010101010001100;
        rom[278] = 24'b000011101001001000101011;
        rom[279] = 24'b000011011101011000011000;
        rom[280] = 24'b000010011101010110001110;
        rom[281] = 24'b000001110010111110100111;
        rom[282] = 24'b000010010110001001011000;
        rom[283] = 24'b000011010101001110110010;
        rom[284] = 24'b000011110101101001111001;
        rom[285] = 24'b000011000100011101100000;
        rom[286] = 24'b000010000101111010001000;
        rom[287] = 24'b000001111010111001111111;
        rom[288] = 24'b000010110010001110010000;
        rom[289] = 24'b000011110000110111010000;
        rom[290] = 24'b000011101101001011110111;
        rom[291] = 24'b000010100111010011101111;
        rom[292] = 24'b000001110110000111010110;
        rom[293] = 24'b000010001010010101001101;
        rom[294] = 24'b000011010000101111011000;
        rom[295] = 24'b000011110011111010001000;
        rom[296] = 24'b000011001110011011000001;
        rom[297] = 24'b000010010011010001010111;
        rom[298] = 24'b000010001001111101010100;
        rom[299] = 24'b000010111011100011010011;
        rom[300] = 24'b000011110101101110101010;
        rom[301] = 24'b000011110101010011110100;
        rom[302] = 24'b000011000010011110101011;
        rom[303] = 24'b000010010010000111110110;
        rom[304] = 24'b000010100011011001110111;
        rom[305] = 24'b000011110011000101000110;
        rom[306] = 24'b000100011000110000110000;
        rom[307] = 24'b000011111100110110000110;
        rom[308] = 24'b000010111110010000100111;
        rom[309] = 24'b000010101000000110000110;
        rom[310] = 24'b000011010011100100011011;
        rom[311] = 24'b000100001000110101110100;
        rom[312] = 24'b000100010000100101011010;
        rom[313] = 24'b000011010011111101110011;
        rom[314] = 24'b000010011111111011100100;
        rom[315] = 24'b000010101110001000000111;
        rom[316] = 24'b000011101011101110000001;
        rom[317] = 24'b000100010001001101001000;
        rom[318] = 24'b000011110000011110100111;
        rom[319] = 24'b000010110001011001001101;
        rom[320] = 24'b000010011111100111100110;
        rom[321] = 24'b000011010000110011111111;
        rom[322] = 24'b000100010001110011100111;
        rom[323] = 24'b000100000110110101100000;
        rom[324] = 24'b000010111011111111001111;
        rom[325] = 24'b000010000100101010111111;
        rom[326] = 24'b000010000101111010001000;
        rom[327] = 24'b000010111111100101000000;
        rom[328] = 24'b000011100010000111111001;
        rom[329] = 24'b000011001001000001100010;
        rom[330] = 24'b000010001001111100000111;
        rom[331] = 24'b000001110000100010010111;
        rom[332] = 24'b000010010110000001011110;
        rom[333] = 24'b000011011000011111111000;
        rom[334] = 24'b000011100001110011111011;
        rom[335] = 24'b000010100110011100111100;
        rom[336] = 24'b000001101001110101010101;
        rom[337] = 24'b000001101111001000101011;
        rom[338] = 24'b000010101011101110110100;
        rom[339] = 24'b000011010111001101001001;
        rom[340] = 24'b000011000101111011001000;
        rom[341] = 24'b000010000000000000111001;
        rom[342] = 24'b000001101000111110110000;
        rom[343] = 24'b000010001001110001111001;
        rom[344] = 24'b000011001101001111111000;
        rom[345] = 24'b000011100101110110101001;
        rom[346] = 24'b000010101001010010100100;
        rom[347] = 24'b000001100111110011111011;
        rom[348] = 24'b000001101100010001100101;
        rom[349] = 24'b000010101011010101011100;
        rom[350] = 24'b000011100001110011111011;
        rom[351] = 24'b000011010001001011001000;
        rom[352] = 24'b000010000111010111111110;
        rom[353] = 24'b000001011000000111110111;
        rom[354] = 24'b000001111000110110011000;
        rom[355] = 24'b000010110000100111000010;
        rom[356] = 24'b000010110011101111001001;
        rom[357] = 24'b000001111101101010010000;
        rom[358] = 24'b000000110000011101011000;
        rom[359] = 24'b000000010110110011101111;
        rom[360] = 24'b000001000001111010110000;
        rom[361] = 24'b000010000111111000100000;
        rom[362] = 24'b000010101011010001000111;
        rom[363] = 24'b000010100100110111011111;
        rom[364] = 24'b000010111100111010100110;
        rom[365] = 24'b000100011100110100001101;
        rom[366] = 24'b000111011000011010011000;
        rom[367] = 24'b001001110011001101011000;
        rom[368] = 24'b001010111011100101100001;
        rom[369] = 24'b001011000111001111000111;
        rom[370] = 24'b001011011000110001110100;
        rom[371] = 24'b001011111011101110010011;
        rom[372] = 24'b001011101100101010001010;
        rom[373] = 24'b001001101000011001110100;
        rom[374] = 24'b000110001101000111011011;
        rom[375] = 24'b000011010110011110110110;
        rom[376] = 24'b000010011100000101000111;
        rom[377] = 24'b000010100010100000110110;
        rom[378] = 24'b000010101000011101010000;
        rom[379] = 24'b000001111001000000100110;
        rom[380] = 24'b000001000001101111110111;
        rom[381] = 24'b000000111100101011000110;
        rom[382] = 24'b000001111110000111101011;
        rom[383] = 24'b000010111010101101110100;
        rom[384] = 24'b000011000000000001001010;
        rom[385] = 24'b000010000011011001100011;
        rom[386] = 24'b000001010100001111110100;
        rom[387] = 24'b000001100010011100010111;
        rom[388] = 24'b000010100010011110100001;
        rom[389] = 24'b000011000011000101001000;
        rom[390] = 24'b000010101001101011011000;
        rom[391] = 24'b000001101000001001101101;
        rom[392] = 24'b000001001111000011010110;
        rom[393] = 24'b000010000000001111101111;
        rom[394] = 24'b000010110101000010000111;
        rom[395] = 24'b000010110110010001010000;
        rom[396] = 24'b000001111110111100111111;
        rom[397] = 24'b000001001100100001001111;
        rom[398] = 24'b000001010111100001011000;
        rom[399] = 24'b000010011000100001000000;
        rom[400] = 24'b000010111101100000001001;
        rom[401] = 24'b000010101001010010010010;
        rom[402] = 24'b000001101100101001001000;
        rom[403] = 24'b000001010011001111010111;
        rom[404] = 24'b000001110011110101111110;
        rom[405] = 24'b000010110011111000001000;
        rom[406] = 24'b000010111010101111111011;
        rom[407] = 24'b000010000100010001011100;
        rom[408] = 24'b000001001010000110000101;
        rom[409] = 24'b000001010110101110001011;
        rom[410] = 24'b000010010011010100010100;
        rom[411] = 24'b000011000001001110111001;
        rom[412] = 24'b000010101000101000001000;
        rom[413] = 24'b000001100010101101111001;
        rom[414] = 24'b000001000110110011010000;
        rom[415] = 24'b000001100101001010001001;
        rom[416] = 24'b000010101000101000001000;
        rom[417] = 24'b000010111001111010001001;
        rom[418] = 24'b000010000111000111000100;
        rom[419] = 24'b000001001100111101001011;
        rom[420] = 24'b000001001110111110100101;
        rom[421] = 24'b000010001001001001111100;
        rom[422] = 24'b000010111111101000011011;
        rom[423] = 24'b000010110011111000001000;
        rom[424] = 24'b000001101100100001001110;
        rom[425] = 24'b000001000010001001100111;
        rom[426] = 24'b000001101010001100111000;
        rom[427] = 24'b000010101011101110100010;
        rom[428] = 24'b000011000111010001001001;
        rom[429] = 24'b000010011010111101010000;
        rom[430] = 24'b000001010000001100101000;
        rom[431] = 24'b000001001010000100111111;
        rom[432] = 24'b000010000110010001110000;
        rom[433] = 24'b000011000000000010010000;
        rom[434] = 24'b000010111110110011000111;
        rom[435] = 24'b000001111000111010111111;
        rom[436] = 24'b000001001010001010110110;
        rom[437] = 24'b000001011011111100011101;
        rom[438] = 24'b000010100010010110101000;
        rom[439] = 24'b000011000101100001011000;
        rom[440] = 24'b000010011101100110000001;
        rom[441] = 24'b000001100000000000000111;
        rom[442] = 24'b000001001000000010100100;
        rom[443] = 24'b000001110111001100010011;
        rom[444] = 24'b000010110001010111101010;
        rom[445] = 24'b000010110101110101010100;
        rom[446] = 24'b000001111011101011011011;
        rom[447] = 24'b000001000110011100000110;
        rom[448] = 24'b000001010101010001110111;
        rom[449] = 24'b000010010011110111010110;
        rom[450] = 24'b000010110111000110110000;
        rom[451] = 24'b000010011000101111110110;
        rom[452] = 24'b000001010101010001110111;
        rom[453] = 24'b000000111100101011000110;
        rom[454] = 24'b000001101111011110001011;
        rom[455] = 24'b000010100100101111100100;
        rom[456] = 24'b000010101010000010111010;
        rom[457] = 24'b000001101111110111100011;
        rom[458] = 24'b000001000000101101110100;
        rom[459] = 24'b000001001010000001110111;
        rom[460] = 24'b000010000000010011000001;
        rom[461] = 24'b000010100101110010001000;
        rom[462] = 24'b000010001001111100000111;
        rom[463] = 24'b000001001111101111001101;
        rom[464] = 24'b000000110001110000010110;
        rom[465] = 24'b000001011011100111111111;
        rom[466] = 24'b000010010111101111000111;
        rom[467] = 24'b000010011000111110010000;
        rom[468] = 24'b000001100110100010011111;
        rom[469] = 24'b000000110001101010011111;
        rom[470] = 24'b000000111100101010101000;
        rom[471] = 24'b000001111000110001110000;
        rom[472] = 24'b000010011101110000111001;
        rom[473] = 24'b000010000010001110010010;
        rom[474] = 24'b000001001000000001011000;
        rom[475] = 24'b000000101110100111100111;
        rom[476] = 24'b000001011000111111001110;
        rom[477] = 24'b000010011011011101101000;
        rom[478] = 24'b000010101100000110011011;
        rom[479] = 24'b000001110101100111111100;
        rom[480] = 24'b000001001010000110000101;
        rom[481] = 24'b000001010100010001111011;
        rom[482] = 24'b000010011101000101010100;
        rom[483] = 24'b000011001111111000011001;
        rom[484] = 24'b000010111110100110011000;
        rom[485] = 24'b000001111011001000011001;
        rom[486] = 24'b000001100100000110010000;
        rom[487] = 24'b000010001110101010011001;
        rom[488] = 24'b000011010100100100101000;
        rom[489] = 24'b000011100101110110101001;
        rom[490] = 24'b000010110000100111010100;
        rom[491] = 24'b000001110100000001001011;
        rom[492] = 24'b000001110110000010100101;
        rom[493] = 24'b000010110101000110011100;
        rom[494] = 24'b000011101110000001001011;
        rom[495] = 24'b000011011111110100101000;
        rom[496] = 24'b000010010110000001011110;
        rom[497] = 24'b000001101110000110000111;
        rom[498] = 24'b000010001110110100101000;
        rom[499] = 24'b000011010101001110110010;
        rom[500] = 24'b000011101110010101001001;
        rom[501] = 24'b000011000110111001110000;
        rom[502] = 24'b000001111100001001001000;
        rom[503] = 24'b000001101110101100101111;
        rom[504] = 24'b000010110010001110001111;
        rom[505] = 24'b000011100111000110010000;
        rom[506] = 24'b000011100011011010110111;
        rom[507] = 24'b000010100100110111011111;
        rom[508] = 24'b000001101110110010100110;
        rom[509] = 24'b000010000101011100101101;
        rom[510] = 24'b000011001110010011001000;
        rom[511] = 24'b000011101111000001101000;
        rom[512] = 24'b000011000010001101110001;
        rom[513] = 24'b000010000111000100000111;
        rom[514] = 24'b000001110011111111000100;
        rom[515] = 24'b000010101000000001010011;
        rom[516] = 24'b000011100100101000111010;
        rom[517] = 24'b000011101001000110100100;
        rom[518] = 24'b000010101110111100101011;
        rom[519] = 24'b000001110111010001000110;
        rom[520] = 24'b000010001000100011000111;
        rom[521] = 24'b000011000100101100010110;
        rom[522] = 24'b000011101010011000000000;
        rom[523] = 24'b000011001110011101010110;
        rom[524] = 24'b000010000110000110110111;
        rom[525] = 24'b000001110010011000100110;
        rom[526] = 24'b000010100010101111011011;
        rom[527] = 24'b000011011000000000110100;
        rom[528] = 24'b000011100010001100101010;
        rom[529] = 24'b000010100101100101000011;
        rom[530] = 24'b000001110011111111000100;
        rom[531] = 24'b000001111101010011000111;
        rom[532] = 24'b000010111000011100110001;
        rom[533] = 24'b000011011101111011111000;
        rom[534] = 24'b000011000010000101110111;
        rom[535] = 24'b000010000000100100001101;
        rom[536] = 24'b000001101001111010000110;
        rom[537] = 24'b000010011000101010001111;
        rom[538] = 24'b000011001101011100100111;
        rom[539] = 24'b000011010011100100010000;
        rom[540] = 24'b000010011110101100001111;
        rom[541] = 24'b000001101100010000011111;
        rom[542] = 24'b000001110111010000101000;
        rom[543] = 24'b000010110101110100000000;
        rom[544] = 24'b000011011010110011001001;
        rom[545] = 24'b000011000001101100110010;
        rom[546] = 24'b000010000000001011000111;
        rom[547] = 24'b000001101110000110000111;
        rom[548] = 24'b000010010001001000111110;
        rom[549] = 24'b000011001110101110111000;
        rom[550] = 24'b000011011010011111001011;
        rom[551] = 24'b000010011111001000001100;
        rom[552] = 24'b000001101110101101110101;
        rom[553] = 24'b000001110100000001001011;
        rom[554] = 24'b000010110000100111010100;
        rom[555] = 24'b000011011110100001111001;
        rom[556] = 24'b000011000001000010101000;
        rom[557] = 24'b000001111101100100101001;
        rom[558] = 24'b000001011100110001100000;
        rom[559] = 24'b000010000010011101001001;
        rom[560] = 24'b000011001000010111011000;
        rom[561] = 24'b000011011001101001011001;
        rom[562] = 24'b000010101001010010100100;
        rom[563] = 24'b000001101100101100011011;
        rom[564] = 24'b000001101001110101010101;
        rom[565] = 24'b000010101011010101011100;
        rom[566] = 24'b000011011111010111101011;
        rom[567] = 24'b000011001110101110111000;
        rom[568] = 24'b000010001001110100001110;
        rom[569] = 24'b000001011111011100100111;
        rom[570] = 24'b000001111101101110111000;
        rom[571] = 24'b000011000100001001000010;
        rom[572] = 24'b000011100010000111111001;
        rom[573] = 24'b000010101110011111010000;
        rom[574] = 24'b000001101111111011111000;
        rom[575] = 24'b000001100010011111011111;
        rom[576] = 24'b000010011100010000000000;
        rom[577] = 24'b000011011000011100110000;
        rom[578] = 24'b000011010100110001010111;
        rom[579] = 24'b000010010001010101011111;
        rom[580] = 24'b000001100101000001100110;
        rom[581] = 24'b000001111110000111111101;
        rom[582] = 24'b000011000100100010001000;
        rom[583] = 24'b000011100000011000001000;
        rom[584] = 24'b000010111010111001000001;
        rom[585] = 24'b000001111000011010100111;
        rom[586] = 24'b000001100101010101100100;
        rom[587] = 24'b000010011001010111110011;
        rom[588] = 24'b000011010101111111011010;
        rom[589] = 24'b000011011000000000110100;
        rom[590] = 24'b000010100010101111011011;
        rom[591] = 24'b000001111100001001100110;
        rom[592] = 24'b000010001101011011100111;
        rom[593] = 24'b000011010000111001100110;
        rom[594] = 24'b000011111001000001100000;
        rom[595] = 24'b000011011010101010100110;
        rom[596] = 24'b000010011110100001010111;
        rom[597] = 24'b000010001010110011000110;
        rom[598] = 24'b000010111011001001111011;
        rom[599] = 24'b000011111100101000100100;
        rom[600] = 24'b000100000001111011111010;
        rom[601] = 24'b000011001100101001000011;
        rom[602] = 24'b000010011111111011100100;
        rom[603] = 24'b000010110011000000100111;
        rom[604] = 24'b000011100110110101100001;
        rom[605] = 24'b000100001100010100101000;
        rom[606] = 24'b000011110000011110100111;
        rom[607] = 24'b000010101100100000101101;
        rom[608] = 24'b000010011000010010110110;
        rom[609] = 24'b000010111111101110001111;
        rom[610] = 24'b000011111011110101010111;
        rom[611] = 24'b000011111000001100000000;
        rom[612] = 24'b000011000000110111101111;
        rom[613] = 24'b000010001110011011111111;
        rom[614] = 24'b000010011110010100101000;
        rom[615] = 24'b000011101001000101010000;
        rom[616] = 24'b000100010111110101011001;
        rom[617] = 24'b000011111001110110100010;
        rom[618] = 24'b000010100111001111000111;
        rom[619] = 24'b000010000110100000100111;
        rom[620] = 24'b000010101001100011011110;
        rom[621] = 24'b000011100111001001011000;
        rom[622] = 24'b000011101011100100111011;
        rom[623] = 24'b000010110000001101111100;
        rom[624] = 24'b000001101100010001100101;
        rom[625] = 24'b000001110100000001001011;
        rom[626] = 24'b000010101110001011000100;
        rom[627] = 24'b000011011110100001111001;
        rom[628] = 24'b000011000001000010101000;
        rom[629] = 24'b000001111000101100001001;
        rom[630] = 24'b000001011010010101010000;
        rom[631] = 24'b000010000100111001011001;
        rom[632] = 24'b000011000011011110111000;
        rom[633] = 24'b000011010100110000111001;
        rom[634] = 24'b000010011111100001100100;
        rom[635] = 24'b000001011110000010111011;
        rom[636] = 24'b000001011000101111100101;
        rom[637] = 24'b000010010111110011011100;
        rom[638] = 24'b000011001110010001111011;
        rom[639] = 24'b000011000000000101011000;
        rom[640] = 24'b000001111000101110011110;
        rom[641] = 24'b000001001110010110110111;
        rom[642] = 24'b000001101111000101010111;
        rom[643] = 24'b000010110011000011010010;
        rom[644] = 24'b000011010101111010101001;
        rom[645] = 24'b000010100010010010000000;
        rom[646] = 24'b000001011001111101101000;
        rom[647] = 24'b000001001010000100111111;
        rom[648] = 24'b000001111110111101000000;
        rom[649] = 24'b000010101010000100000000;
        rom[650] = 24'b000010010010110110100111;
        rom[651] = 24'b000001001000000101111111;
        rom[652] = 24'b000000001101001000100110;
        rom[653] = 24'b000000010101001001001101;
        rom[654] = 24'b000001001111010110001000;
        rom[655] = 24'b000010000011100110101000;
        rom[656] = 24'b000010010110010001010001;
        rom[657] = 24'b000010100001111010110111;
        rom[658] = 24'b000011100001110110010100;
        rom[659] = 24'b000101111100011011000011;
        rom[660] = 24'b001001000100001100111010;
        rom[661] = 24'b001011001010000011110100;
        rom[662] = 24'b001011101100101011011011;
        rom[663] = 24'b001011100000111100010110;
        rom[664] = 24'b001010111110111101000111;
        rom[665] = 24'b001001011110110110010110;
        rom[666] = 24'b000110011100100110010000;
        rom[667] = 24'b000011000100101100010110;
        rom[668] = 24'b000000101011110001100111;
        rom[669] = 24'b000000010101100111000110;
        rom[670] = 24'b000001100011010000111011;
        rom[671] = 24'b000010101110100000100100;
        rom[672] = 24'b000010111011001000101010;
        rom[673] = 24'b000010000011011001100011;
        rom[674] = 24'b000001001100111011000100;
        rom[675] = 24'b000001011101100011110111;
        rom[676] = 24'b000010011011001001110001;
        rom[677] = 24'b000010111110001100101000;
        rom[678] = 24'b000010100100110010110111;
        rom[679] = 24'b000001011110011000101101;
        rom[680] = 24'b000001001100100111000110;
        rom[681] = 24'b000001110110011110101111;
        rom[682] = 24'b000010110101000010000111;
        rom[683] = 24'b000010110110010001010000;
        rom[684] = 24'b000010000001011001001111;
        rom[685] = 24'b000001001100100001001111;
        rom[686] = 24'b000001010101000101001000;
        rom[687] = 24'b000010001100010011110000;
        rom[688] = 24'b000010111101100000001001;
        rom[689] = 24'b000010011101000101000010;
        rom[690] = 24'b000001011101111111100111;
        rom[691] = 24'b000001000100100101110111;
        rom[692] = 24'b000001101100100001001110;
        rom[693] = 24'b000010100101001110101000;
        rom[694] = 24'b000010110011011011001011;
        rom[695] = 24'b000001111000000100001100;
        rom[696] = 24'b000001000101001101100101;
        rom[697] = 24'b000001001100111101001011;
        rom[698] = 24'b000010001001100011010100;
        rom[699] = 24'b000010111100010110011001;
        rom[700] = 24'b000010011110110111001000;
        rom[701] = 24'b000001011011011001001001;
        rom[702] = 24'b000000111101000010010000;
        rom[703] = 24'b000001100010101101111001;
        rom[704] = 24'b000010100110001011111000;
        rom[705] = 24'b000010111001111010001001;
        rom[706] = 24'b000010000010001110100100;
        rom[707] = 24'b000001001000000100101011;
        rom[708] = 24'b000001001110111110100101;
        rom[709] = 24'b000010001011100110001100;
        rom[710] = 24'b000010111101001100001011;
        rom[711] = 24'b000010101110111111101000;
        rom[712] = 24'b000001110001011001101110;
        rom[713] = 24'b000000111111101101010111;
        rom[714] = 24'b000001100010111000001000;
        rom[715] = 24'b000010101011101110100010;
        rom[716] = 24'b000010111111111100011001;
        rom[717] = 24'b000010010011101000100000;
        rom[718] = 24'b000001001101110000011000;
        rom[719] = 24'b000001000000010011111111;
        rom[720] = 24'b000001110111101000010000;
        rom[721] = 24'b000010110011110101000000;
        rom[722] = 24'b000010101011010001000111;
        rom[723] = 24'b000001101111001001111111;
        rom[724] = 24'b000000111011100001010110;
        rom[725] = 24'b000001010100100111101101;
        rom[726] = 24'b000010011000100101101000;
        rom[727] = 24'b000010111001010100001000;
        rom[728] = 24'b000010011000101101100001;
        rom[729] = 24'b000001011000101011010111;
        rom[730] = 24'b000001000101100110010100;
        rom[731] = 24'b000001110010010011110011;
        rom[732] = 24'b000010110011110011111010;
        rom[733] = 24'b000010110011011001000100;
        rom[734] = 24'b000001111011101011011011;
        rom[735] = 24'b000001001000111000010110;
        rom[736] = 24'b000001011100100110100111;
        rom[737] = 24'b000010011011001100000110;
        rom[738] = 24'b000011001000001100100000;
        rom[739] = 24'b000010011101101000010110;
        rom[740] = 24'b000001100001011111000111;
        rom[741] = 24'b000001001101110000110110;
        rom[742] = 24'b000001111001001111001011;
        rom[743] = 24'b000010101110100000100100;
        rom[744] = 24'b000010110110010000001010;
        rom[745] = 24'b000001111100000100110011;
        rom[746] = 24'b000001000101100110010100;
        rom[747] = 24'b000001010001010110100111;
        rom[748] = 24'b000010001110111100100001;
        rom[749] = 24'b000010110110110111111000;
        rom[750] = 24'b000010010110001001010111;
        rom[751] = 24'b000001011001100000001101;
        rom[752] = 24'b000001000000011001110110;
        rom[753] = 24'b000001101111001001111111;
        rom[754] = 24'b000010100001100000000111;
        rom[755] = 24'b000010101100100000010000;
        rom[756] = 24'b000001110010101111101111;
        rom[757] = 24'b000001000010110000001111;
        rom[758] = 24'b000001001011010100001000;
        rom[759] = 24'b000010001001110111100000;
        rom[760] = 24'b000010110110001011011001;
        rom[761] = 24'b000010011010101000110010;
        rom[762] = 24'b000001011001000111000111;
        rom[763] = 24'b000000111111101101010111;
        rom[764] = 24'b000001110001011001101110;
        rom[765] = 24'b000010110001011011111000;
        rom[766] = 24'b000011000010000100101011;
        rom[767] = 24'b000010010101010111001100;
        rom[768] = 24'b000001100010100000100101;
        rom[769] = 24'b000001101111001000101011;
        rom[770] = 24'b000010101110001011000100;
        rom[771] = 24'b000011100000111110001001;
        rom[772] = 24'b000011001010110011101000;
        rom[773] = 24'b000010001001110001111001;
        rom[774] = 24'b000001101011011011000000;
        rom[775] = 24'b000010010001000110101001;
        rom[776] = 24'b000011011001011101001000;
        rom[777] = 24'b000011101101001011011001;
        rom[778] = 24'b000010110111111100000100;
        rom[779] = 24'b000001111101110010001011;
        rom[780] = 24'b000001111101010111010101;
        rom[781] = 24'b000010111001111110111100;
        rom[782] = 24'b000011101110000001001011;
        rom[783] = 24'b000011011111110100101000;
        rom[784] = 24'b000010011010111001111110;
        rom[785] = 24'b000001110010111110100111;
        rom[786] = 24'b000010010001010000111000;
        rom[787] = 24'b000011010000010110010010;
        rom[788] = 24'b000011110000110001011001;
        rom[789] = 24'b000011000010000001010000;
        rom[790] = 24'b000001111110100101011000;
        rom[791] = 24'b000001110011100101001111;
        rom[792] = 24'b000010101000011101010000;
        rom[793] = 24'b000011100111000110010000;
        rom[794] = 24'b000011100000111110100111;
        rom[795] = 24'b000010100010011011001111;
        rom[796] = 24'b000001101110110010100110;
        rom[797] = 24'b000010000101011100101101;
        rom[798] = 24'b000011010000101111010111;
        rom[799] = 24'b000011101100100101011000;
        rom[800] = 24'b000011001011111110110001;
        rom[801] = 24'b000010000100100111110111;
        rom[802] = 24'b000001101111000110100100;
        rom[803] = 24'b000010100000101100100011;
        rom[804] = 24'b000011011111110000011010;
        rom[805] = 24'b000011011100111001010100;
        rom[806] = 24'b000010100000010011001011;
        rom[807] = 24'b000001101101100000000110;
        rom[808] = 24'b000001110101000001000111;
        rom[809] = 24'b000010110110000010110110;
        rom[810] = 24'b000011011110001010110000;
        rom[811] = 24'b000010111101010111100110;
        rom[812] = 24'b000001111110110010000111;
        rom[813] = 24'b000001101000100111100110;
        rom[814] = 24'b000010010110100010001011;
        rom[815] = 24'b000011001001010111010100;
        rom[816] = 24'b000011010001000110111010;
        rom[817] = 24'b000010010110111011100011;
        rom[818] = 24'b000001100000011101000100;
        rom[819] = 24'b000001101100001101010111;
        rom[820] = 24'b000010101110101011110001;
        rom[821] = 24'b000011010001101110101000;
        rom[822] = 24'b000010111000010100110111;
        rom[823] = 24'b000001111001001111011101;
        rom[824] = 24'b000001100101000001100110;
        rom[825] = 24'b000010001010000000101111;
        rom[826] = 24'b000011001011000000010111;
        rom[827] = 24'b000011001100001111100000;
        rom[828] = 24'b000010010100111011010000;
        rom[829] = 24'b000001100100111011101111;
        rom[830] = 24'b000001101011000011011000;
        rom[831] = 24'b000010101100000011000000;
        rom[832] = 24'b000011001110100101111001;
        rom[833] = 24'b000010110000100111000010;
        rom[834] = 24'b000001110011111101110111;
        rom[835] = 24'b000001011010100100000111;
        rom[836] = 24'b000010000000000011001110;
        rom[837] = 24'b000011000010100001101000;
        rom[838] = 24'b000011001110010001111011;
        rom[839] = 24'b000010010010111010111100;
        rom[840] = 24'b000001011101101000000101;
        rom[841] = 24'b000001100010111011011011;
        rom[842] = 24'b000010100110110110010100;
        rom[843] = 24'b000011010111001101001001;
        rom[844] = 24'b000011000011011110111000;
        rom[845] = 24'b000001111000101100001001;
        rom[846] = 24'b000001010111111001000000;
        rom[847] = 24'b000010000100111001011001;
        rom[848] = 24'b000011000101111011001000;
        rom[849] = 24'b000011011100000101101001;
        rom[850] = 24'b000010100100011010000100;
        rom[851] = 24'b000001100010111011011011;
        rom[852] = 24'b000001100010100000100101;
        rom[853] = 24'b000010011111001000001100;
        rom[854] = 24'b000011010011001010011011;
        rom[855] = 24'b000011000100111101111000;
        rom[856] = 24'b000001111011001010101110;
        rom[857] = 24'b000001001110010110110111;
        rom[858] = 24'b000001111011010010101000;
        rom[859] = 24'b000010111010011000000010;
        rom[860] = 24'b000011010101111010101001;
        rom[861] = 24'b000010100111001010100000;
        rom[862] = 24'b000001101000100111001000;
        rom[863] = 24'b000001011011001010101111;
        rom[864] = 24'b000010010111010111100000;
        rom[865] = 24'b000011010110000000100000;
        rom[866] = 24'b000011001000100100000111;
        rom[867] = 24'b000010001110111001001111;
        rom[868] = 24'b000001100010100101010110;
        rom[869] = 24'b000001111011101011101101;
        rom[870] = 24'b000010111111101001101000;
        rom[871] = 24'b000011101100100101011000;
        rom[872] = 24'b000011000111000110010001;
        rom[873] = 24'b000010000111000100000111;
        rom[874] = 24'b000001110110011011010100;
        rom[875] = 24'b000010101100111001110011;
        rom[876] = 24'b000011101110011001111010;
        rom[877] = 24'b000011101101111111000100;
        rom[878] = 24'b000010110110010001011011;
        rom[879] = 24'b000010000011011110010110;
        rom[880] = 24'b000010010111001100100111;
        rom[881] = 24'b000011011010101010100110;
        rom[882] = 24'b000100000010110010100000;
        rom[883] = 24'b000011100100011011100110;
        rom[884] = 24'b000010101000010010010111;
        rom[885] = 24'b000010001101001111010110;
        rom[886] = 24'b000010111011001001111011;
        rom[887] = 24'b000011110010110111100100;
        rom[888] = 24'b000011110011010010011010;
        rom[889] = 24'b000011000000011011110011;
        rom[890] = 24'b000010001001111101010100;
        rom[891] = 24'b000010010101101101100111;
        rom[892] = 24'b000011010011010011100001;
        rom[893] = 24'b000011111101101011001000;
        rom[894] = 24'b000011011100111100100111;
        rom[895] = 24'b000010011101110111001101;
        rom[896] = 24'b000010001001101001010110;
        rom[897] = 24'b000010111010110101101111;
        rom[898] = 24'b000100000000101101110111;
        rom[899] = 24'b000011111111100000110000;
        rom[900] = 24'b000010111110011011011111;
        rom[901] = 24'b000001111000011101101111;
        rom[902] = 24'b000010000001000001101000;
        rom[903] = 24'b000010101110011111010000;
        rom[904] = 24'b000011010011011110011001;
        rom[905] = 24'b000010110000100111000010;
        rom[906] = 24'b000001101100101001001000;
        rom[907] = 24'b000001010000110011000111;
        rom[908] = 24'b000001111101100110111110;
        rom[909] = 24'b000010111011001100111000;
        rom[910] = 24'b000011000100100000111011;
        rom[911] = 24'b000010001110000010011100;
        rom[912] = 24'b000001010001011010110101;
        rom[913] = 24'b000001011001001010011011;
        rom[914] = 24'b000010010101110000100100;
        rom[915] = 24'b000011000110000111011001;
        rom[916] = 24'b000010101101100000101000;
        rom[917] = 24'b000001100111100110011001;
        rom[918] = 24'b000001000110110011010000;
        rom[919] = 24'b000001110110001111111001;
        rom[920] = 24'b000010110111010001101000;
        rom[921] = 24'b000011000011101011001001;
        rom[922] = 24'b000010010000111000000100;
        rom[923] = 24'b000001001010100000111011;
        rom[924] = 24'b000001001100100010010101;
        rom[925] = 24'b000010001001001001111100;
        rom[926] = 24'b000011000010000100101011;
        rom[927] = 24'b000010101100100011011000;
        rom[928] = 24'b000001100010110000001110;
        rom[929] = 24'b000000101001101111000111;
        rom[930] = 24'b000001000000101100101000;
        rom[931] = 24'b000001110011100100110010;
        rom[932] = 24'b000010001010001110111001;
        rom[933] = 24'b000001010110100110010000;
        rom[934] = 24'b000000010000101110001000;
        rom[935] = 24'b111111101010110111001111;
        rom[936] = 24'b000000001100001101010000;
        rom[937] = 24'b000001001010110110010000;
        rom[938] = 24'b000001011101001001000111;
        rom[939] = 24'b000001000101101001101111;
        rom[940] = 24'b000001001111000011010110;
        rom[941] = 24'b000010100000010011011101;
        rom[942] = 24'b000100101101100000111000;
        rom[943] = 24'b000110101111111001011000;
        rom[944] = 24'b001000010000101100000001;
        rom[945] = 24'b001001010010000011000111;
        rom[946] = 24'b001010011001010011010100;
        rom[947] = 24'b001011100101110000000011;
        rom[948] = 24'b001011110011111110111010;
        rom[949] = 24'b001001100001000101000100;
        rom[950] = 24'b000101011100010010011011;
        rom[951] = 24'b000001110111010001000110;
        rom[952] = 24'b000000101011110001100111;
        rom[953] = 24'b000001100011000010010110;
        rom[954] = 24'b000010011100010000000000;
        rom[955] = 24'b000010011000101111110110;
        rom[956] = 24'b000001100001011111000111;
        rom[957] = 24'b000001001101110000110110;
        rom[958] = 24'b000001111001001111001011;
        rom[959] = 24'b000010110000111100110100;
        rom[960] = 24'b000010110110010000001010;
        rom[961] = 24'b000010000101110101110011;
        rom[962] = 24'b000001001111010111010100;
        rom[963] = 24'b000001011011000111100111;
        rom[964] = 24'b000010010110010001010001;
        rom[965] = 24'b000010111011110000011000;
        rom[966] = 24'b000010011111111010010111;
        rom[967] = 24'b000001100000110100111101;
        rom[968] = 24'b000001001100100111000110;
        rom[969] = 24'b000001110110011110101111;
        rom[970] = 24'b000010101101101101010111;
        rom[971] = 24'b000010110011110101000000;
        rom[972] = 24'b000001111110111101000000;
        rom[973] = 24'b000001001110111101011111;
        rom[974] = 24'b000001010010101000111000;
        rom[975] = 24'b000010001110110000000000;
        rom[976] = 24'b000010111101100000001001;
        rom[977] = 24'b000010100100011001110010;
        rom[978] = 24'b000001100000011011110111;
        rom[979] = 24'b000001001011111010100111;
        rom[980] = 24'b000001110110010010001110;
        rom[981] = 24'b000010110011111000001000;
        rom[982] = 24'b000010111111101000011011;
        rom[983] = 24'b000010001001001001111100;
        rom[984] = 24'b000001001110111110100101;
        rom[985] = 24'b000001010001110101101011;
        rom[986] = 24'b000010010000111000000100;
        rom[987] = 24'b000011000001001110111001;
        rom[988] = 24'b000010101000101000001000;
        rom[989] = 24'b000001100111100110011001;
        rom[990] = 24'b000001000110110011010000;
        rom[991] = 24'b000001101100011110111001;
        rom[992] = 24'b000010110010011001001000;
        rom[993] = 24'b000011001010111111111001;
        rom[994] = 24'b000010010101110000100100;
        rom[995] = 24'b000001010100010001111011;
        rom[996] = 24'b000001010011110111000101;
        rom[997] = 24'b000010010000011110101100;
        rom[998] = 24'b000011001001011001011011;
        rom[999] = 24'b000010110110010100011000;
        rom[1000] = 24'b000001110001011001101110;
        rom[1001] = 24'b000001001001011110010111;
        rom[1002] = 24'b000001101100101001001000;
        rom[1003] = 24'b000010110011000011010010;
        rom[1004] = 24'b000011001100001001101001;
        rom[1005] = 24'b000010011010111101010000;
        rom[1006] = 24'b000001010111100001011000;
        rom[1007] = 24'b000001010001011001101111;
        rom[1008] = 24'b000010001000101101111111;
        rom[1009] = 24'b000011001100001111100000;
        rom[1010] = 24'b000010111110110011000111;
        rom[1011] = 24'b000001111011010111001111;
        rom[1012] = 24'b000001001010001010110110;
        rom[1013] = 24'b000001101010100101111101;
        rom[1014] = 24'b000010101001101011011000;
        rom[1015] = 24'b000011001100110110001000;
        rom[1016] = 24'b000010100010011110100001;
        rom[1017] = 24'b000001011101100011110111;
        rom[1018] = 24'b000001010100001111110100;
        rom[1019] = 24'b000010001010101110010011;
        rom[1020] = 24'b000011000100111001101010;
        rom[1021] = 24'b000011000010000010100100;
        rom[1022] = 24'b000010000101011100011011;
        rom[1023] = 24'b000001010010101001010110;
        rom[1024] = 24'b000001100001011111000111;
        rom[1025] = 24'b000010100010100000110110;
        rom[1026] = 24'b000011010001111101100000;
        rom[1027] = 24'b000010101100010001110110;
        rom[1028] = 24'b000001101000110011110111;
        rom[1029] = 24'b000001010000001101000110;
        rom[1030] = 24'b000001111110000111101011;
        rom[1031] = 24'b000010111010101101110100;
        rom[1032] = 24'b000011000100111001101010;
        rom[1033] = 24'b000010001111100110110011;
        rom[1034] = 24'b000001010001110011100100;
        rom[1035] = 24'b000001100010011100010111;
        rom[1036] = 24'b000010011101100110000001;
        rom[1037] = 24'b000011001100110110001000;
        rom[1038] = 24'b000010101110100011110111;
        rom[1039] = 24'b000001110001111010101101;
        rom[1040] = 24'b000001010110011000000110;
        rom[1041] = 24'b000001111011010111001111;
        rom[1042] = 24'b000010110101000010000111;
        rom[1043] = 24'b000011000010011110100000;
        rom[1044] = 24'b000010001011001010001111;
        rom[1045] = 24'b000001011011001010101111;
        rom[1046] = 24'b000001100110001010111000;
        rom[1047] = 24'b000010100010010010000000;
        rom[1048] = 24'b000011001100001001101001;
        rom[1049] = 24'b000010111111010000100010;
        rom[1050] = 24'b000010000101000011100111;
        rom[1051] = 24'b000001101110000110000111;
        rom[1052] = 24'b000010011000011101101110;
        rom[1053] = 24'b000011010110000011101000;
        rom[1054] = 24'b000011100001110011111011;
        rom[1055] = 24'b000010110010101010001100;
        rom[1056] = 24'b000010000010001111110101;
        rom[1057] = 24'b000010001001111111011011;
        rom[1058] = 24'b000010111111010000110100;
        rom[1059] = 24'b000011110010000011111001;
        rom[1060] = 24'b000011100011001110001000;
        rom[1061] = 24'b000010100010001100011001;
        rom[1062] = 24'b000010000001011001010000;
        rom[1063] = 24'b000010101001100001001001;
        rom[1064] = 24'b000011100101101010011000;
        rom[1065] = 24'b000011110100100000001001;
        rom[1066] = 24'b000011000001101101000100;
        rom[1067] = 24'b000010000101000110111011;
        rom[1068] = 24'b000010000100101100000101;
        rom[1069] = 24'b000011000011101111111100;
        rom[1070] = 24'b000011110010111001101011;
        rom[1071] = 24'b000011100010010000111000;
        rom[1072] = 24'b000010011010111001111110;
        rom[1073] = 24'b000001111010010011010111;
        rom[1074] = 24'b000010011101011110001000;
        rom[1075] = 24'b000011100001011100000010;
        rom[1076] = 24'b000011111100111110101001;
        rom[1077] = 24'b000011000110111001110000;
        rom[1078] = 24'b000010000011011101111000;
        rom[1079] = 24'b000001111101010110001111;
        rom[1080] = 24'b000010110111000110110000;
        rom[1081] = 24'b000011101110011011000000;
        rom[1082] = 24'b000011101010101111100111;
        rom[1083] = 24'b000010100100110111011111;
        rom[1084] = 24'b000001110110000111010110;
        rom[1085] = 24'b000010010001101001111101;
        rom[1086] = 24'b000011010101100111110111;
        rom[1087] = 24'b000011110001011101111000;
        rom[1088] = 24'b000011000111000110010001;
        rom[1089] = 24'b000010000010001011100111;
        rom[1090] = 24'b000001110110011011010100;
        rom[1091] = 24'b000010101000000001010011;
        rom[1092] = 24'b000011101011111101101010;
        rom[1093] = 24'b000011100110101010010100;
        rom[1094] = 24'b000010100101001011101011;
        rom[1095] = 24'b000001101011000011110110;
        rom[1096] = 24'b000001111001111001100111;
        rom[1097] = 24'b000010111111110011110110;
        rom[1098] = 24'b000011100111111011110000;
        rom[1099] = 24'b000011000100101100010110;
        rom[1100] = 24'b000010000110000110110111;
        rom[1101] = 24'b000001101101100000000110;
        rom[1102] = 24'b000010011000111110011011;
        rom[1103] = 24'b000011011000000000110100;
        rom[1104] = 24'b000011100010001100101010;
        rom[1105] = 24'b000010100101100101000011;
        rom[1106] = 24'b000001110001100010110100;
        rom[1107] = 24'b000001111010110110110111;
        rom[1108] = 24'b000010110011100100010001;
        rom[1109] = 24'b000011011101111011111000;
        rom[1110] = 24'b000011000010000101111000;
        rom[1111] = 24'b000010000011000000011101;
        rom[1112] = 24'b000001100111011101110110;
        rom[1113] = 24'b000010001110111001001111;
        rom[1114] = 24'b000011001011000000010111;
        rom[1115] = 24'b000011010110000000100000;
        rom[1116] = 24'b000010100001001000011111;
        rom[1117] = 24'b000001101100010000011111;
        rom[1118] = 24'b000001110100110100011000;
        rom[1119] = 24'b000010110101110100000000;
        rom[1120] = 24'b000011011111101011101001;
        rom[1121] = 24'b000011000100001001000010;
        rom[1122] = 24'b000010000101000011100111;
        rom[1123] = 24'b000001101110000110000111;
        rom[1124] = 24'b000010001100010000011110;
        rom[1125] = 24'b000011001100010010101000;
        rom[1126] = 24'b000011010101100110101011;
        rom[1127] = 24'b000010011010001111101100;
        rom[1128] = 24'b000001100010100000100101;
        rom[1129] = 24'b000001101100101100011011;
        rom[1130] = 24'b000010101001010010100100;
        rom[1131] = 24'b000011010111001101001001;
        rom[1132] = 24'b000011000011011110111000;
        rom[1133] = 24'b000010000010011101001001;
        rom[1134] = 24'b000001100100000110010000;
        rom[1135] = 24'b000010000111010101101001;
        rom[1136] = 24'b000011000101111011001000;
        rom[1137] = 24'b000011011001101001011001;
        rom[1138] = 24'b000010011000001100110100;
        rom[1139] = 24'b000001100101010111101011;
        rom[1140] = 24'b000001100010100000100101;
        rom[1141] = 24'b000010100100000000101100;
        rom[1142] = 24'b000011011000000010111011;
        rom[1143] = 24'b000011000111011010001000;
        rom[1144] = 24'b000010000100111011101110;
        rom[1145] = 24'b000001100001111000110111;
        rom[1146] = 24'b000010000111011111111000;
        rom[1147] = 24'b000011001001000001100010;
        rom[1148] = 24'b000011011111101011101001;
        rom[1149] = 24'b000010110011010111110000;
        rom[1150] = 24'b000001110010011000001000;
        rom[1151] = 24'b000001101110101100101111;
        rom[1152] = 24'b000010101010111001100000;
        rom[1153] = 24'b000011110000110111010000;
        rom[1154] = 24'b000011101000010011010111;
        rom[1155] = 24'b000010100100110111011111;
        rom[1156] = 24'b000001110110000111010110;
        rom[1157] = 24'b000010011000111110101101;
        rom[1158] = 24'b000011011100111100100111;
        rom[1159] = 24'b000011111101101011001000;
        rom[1160] = 24'b000011010011010011100001;
        rom[1161] = 24'b000010010101101101100111;
        rom[1162] = 24'b000010001001111101010100;
        rom[1163] = 24'b000011000000011011110011;
        rom[1164] = 24'b000100000001111011111010;
        rom[1165] = 24'b000100001000110101110100;
        rom[1166] = 24'b000011000100111010111011;
        rom[1167] = 24'b000010010111000000010110;
        rom[1168] = 24'b000010100011011001110111;
        rom[1169] = 24'b000011100100011011100110;
        rom[1170] = 24'b000100001100100011100000;
        rom[1171] = 24'b000011101110001100100110;
        rom[1172] = 24'b000010100011011001110111;
        rom[1173] = 24'b000010001010110011000110;
        rom[1174] = 24'b000010111101100110001011;
        rom[1175] = 24'b000011111100101000100100;
        rom[1176] = 24'b000011111000001010111010;
        rom[1177] = 24'b000011000000011011110011;
        rom[1178] = 24'b000010000101000100110100;
        rom[1179] = 24'b000010011111011110100111;
        rom[1180] = 24'b000011100001111101000001;
        rom[1181] = 24'b000100001100010100101000;
        rom[1182] = 24'b000011100100010001010111;
        rom[1183] = 24'b000010011011011010111101;
        rom[1184] = 24'b000001111000100011100110;
        rom[1185] = 24'b000010011101100010101111;
        rom[1186] = 24'b000011010111001101100111;
        rom[1187] = 24'b000011011010111001000000;
        rom[1188] = 24'b000010011110101100001111;
        rom[1189] = 24'b000001101110101100101111;
        rom[1190] = 24'b000001110100110100011000;
        rom[1191] = 24'b000010101110011111010000;
        rom[1192] = 24'b000011010011011110011001;
        rom[1193] = 24'b000010111111010000100010;
        rom[1194] = 24'b000010000010100111010111;
        rom[1195] = 24'b000001100110110001010111;
        rom[1196] = 24'b000010001001110100001110;
        rom[1197] = 24'b000011000010100001101000;
        rom[1198] = 24'b000011001110010001111011;
        rom[1199] = 24'b000010010101010111001100;
        rom[1200] = 24'b000001011101101000000101;
        rom[1201] = 24'b000001100010111011011011;
        rom[1202] = 24'b000010011111100001100100;
        rom[1203] = 24'b000011001000100011101001;
        rom[1204] = 24'b000010110111010001101000;
        rom[1205] = 24'b000001110110001111111001;
        rom[1206] = 24'b000001010111111001000000;
        rom[1207] = 24'b000001111000101100001001;
        rom[1208] = 24'b000010111110100110011000;
        rom[1209] = 24'b000011001101011100001001;
        rom[1210] = 24'b000010011000001100110100;
        rom[1211] = 24'b000001100010111011011011;
        rom[1212] = 24'b000001100010100000100101;
        rom[1213] = 24'b000010100001100100011100;
        rom[1214] = 24'b000011010011001010011011;
        rom[1215] = 24'b000010111101101001001000;
        rom[1216] = 24'b000001110110010010001110;
        rom[1217] = 24'b000001001001011110010111;
        rom[1218] = 24'b000001010110101010111000;
        rom[1219] = 24'b000010010000110111110010;
        rom[1220] = 24'b000010010110011100001001;
        rom[1221] = 24'b000001011011011110110000;
        rom[1222] = 24'b000000000100100000111000;
        rom[1223] = 24'b000000000000110101011111;
        rom[1224] = 24'b000001011111001101110000;
        rom[1225] = 24'b000011010001001000000000;
        rom[1226] = 24'b000100001010011110110111;
        rom[1227] = 24'b000100011100011111101111;
        rom[1228] = 24'b000101100101010111110110;
        rom[1229] = 24'b001000001100000100101101;
        rom[1230] = 24'b001010111101111001111000;
        rom[1231] = 24'b001100010100010101111000;
        rom[1232] = 24'b001011011000111000100001;
        rom[1233] = 24'b001000100001001110000111;
        rom[1234] = 24'b000101010100100110000100;
        rom[1235] = 24'b000011100000001011000011;
        rom[1236] = 24'b000010101110111011011010;
        rom[1237] = 24'b000010000101000000010100;
        rom[1238] = 24'b000001010010001011001011;
        rom[1239] = 24'b000000110000011101110110;
        rom[1240] = 24'b000001010111101110000111;
        rom[1241] = 24'b000010011101101000010110;
        rom[1242] = 24'b000011000101110000010000;
        rom[1243] = 24'b000010100010100000110110;
        rom[1244] = 24'b000001011100100110100111;
        rom[1245] = 24'b000001000110011100000110;
        rom[1246] = 24'b000001101101000001111011;
        rom[1247] = 24'b000010101001101000000100;
        rom[1248] = 24'b000010110110010000001010;
        rom[1249] = 24'b000010000000111101010011;
        rom[1250] = 24'b000001001000000010100100;
        rom[1251] = 24'b000001010110001111000111;
        rom[1252] = 24'b000010010001011000110001;
        rom[1253] = 24'b000010111110001100101000;
        rom[1254] = 24'b000010101001101011010111;
        rom[1255] = 24'b000001100101101101011101;
        rom[1256] = 24'b000001001010001010110110;
        rom[1257] = 24'b000001110110011110101111;
        rom[1258] = 24'b000010110101000010000111;
        rom[1259] = 24'b000010111101100110000000;
        rom[1260] = 24'b000010001011001010010000;
        rom[1261] = 24'b000001010001011001101111;
        rom[1262] = 24'b000001011001111101101000;
        rom[1263] = 24'b000010010011101000100000;
        rom[1264] = 24'b000010110011101111001001;
        rom[1265] = 24'b000010100001111101100010;
        rom[1266] = 24'b000001100101010100010111;
        rom[1267] = 24'b000001001001011110010111;
        rom[1268] = 24'b000001101110111101011110;
        rom[1269] = 24'b000010101100100011011000;
        rom[1270] = 24'b000010110000111110111011;
        rom[1271] = 24'b000010000001110101001100;
        rom[1272] = 24'b000001001100100010010101;
        rom[1273] = 24'b000001001111011001011011;
        rom[1274] = 24'b000010001011111111100100;
        rom[1275] = 24'b000010111001111010001001;
        rom[1276] = 24'b000010100011101111101000;
        rom[1277] = 24'b000001100111100110011001;
        rom[1278] = 24'b000000111101000010010000;
        rom[1279] = 24'b000001100111100110011001;
        rom[1280] = 24'b000010100110001011111000;
        rom[1281] = 24'b000010111001111010001001;
        rom[1282] = 24'b000010000100101010110100;
        rom[1283] = 24'b000001001010100000111011;
        rom[1284] = 24'b000001001100100010010101;
        rom[1285] = 24'b000010001011100110001100;
        rom[1286] = 24'b000010111111101000011011;
        rom[1287] = 24'b000010110001011011111000;
        rom[1288] = 24'b000001101110111101011110;
        rom[1289] = 24'b000001001001011110010111;
        rom[1290] = 24'b000001100111110000101000;
        rom[1291] = 24'b000010100100011001110010;
        rom[1292] = 24'b000010111101100000001001;
        rom[1293] = 24'b000010001001110111100000;
        rom[1294] = 24'b000001000011111111011000;
        rom[1295] = 24'b000001000101001100011111;
        rom[1296] = 24'b000010000001011001010000;
        rom[1297] = 24'b000010111101100110000000;
        rom[1298] = 24'b000010110111011110010111;
        rom[1299] = 24'b000001101100101101101111;
        rom[1300] = 24'b000001000101010010010110;
        rom[1301] = 24'b000001011110011000101101;
        rom[1302] = 24'b000010100010010110101000;
        rom[1303] = 24'b000011000011000101001000;
        rom[1304] = 24'b000010011011001001110001;
        rom[1305] = 24'b000001010110001111000111;
        rom[1306] = 24'b000001000000101101110100;
        rom[1307] = 24'b000001110111001100010011;
        rom[1308] = 24'b000010111000101100011010;
        rom[1309] = 24'b000010111000010001100100;
        rom[1310] = 24'b000001111001001111001011;
        rom[1311] = 24'b000001000110011100000110;
        rom[1312] = 24'b000001010000011001010111;
        rom[1313] = 24'b000010010001011011000110;
        rom[1314] = 24'b000010110100101010100000;
        rom[1315] = 24'b000010010011110111010110;
        rom[1316] = 24'b000001010000011001010111;
        rom[1317] = 24'b000000110000011101110110;
        rom[1318] = 24'b000001100011010000111011;
        rom[1319] = 24'b000010011101011010110100;
        rom[1320] = 24'b000010100111100110101010;
        rom[1321] = 24'b000001101000100010110011;
        rom[1322] = 24'b000000101000010011010100;
        rom[1323] = 24'b000000111101110100100111;
        rom[1324] = 24'b000001111011011010100001;
        rom[1325] = 24'b000010101101000110111000;
        rom[1326] = 24'b000010010001010000110111;
        rom[1327] = 24'b000001010100100111101101;
        rom[1328] = 24'b000000111001000101000110;
        rom[1329] = 24'b000001011110000100001111;
        rom[1330] = 24'b000010011010001011010111;
        rom[1331] = 24'b000010100101001011100000;
        rom[1332] = 24'b000001110101001011111111;
        rom[1333] = 24'b000001000010110000001111;
        rom[1334] = 24'b000001010000001100101000;
        rom[1335] = 24'b000010000111011011010000;
        rom[1336] = 24'b000010110110001011011001;
        rom[1337] = 24'b000010100100011001110010;
        rom[1338] = 24'b000001101111000101010111;
        rom[1339] = 24'b000001010101101011100111;
        rom[1340] = 24'b000010000000000011001110;
        rom[1341] = 24'b000011000000000101011000;
        rom[1342] = 24'b000011001110010001111011;
        rom[1343] = 24'b000010100100000000101100;
        rom[1344] = 24'b000001110001001010000101;
        rom[1345] = 24'b000001111011010101111011;
        rom[1346] = 24'b000010111100110100100100;
        rom[1347] = 24'b000011101101001011011001;
        rom[1348] = 24'b000011010010001000011000;
        rom[1349] = 24'b000010010101111111001001;
        rom[1350] = 24'b000001110010101111110000;
        rom[1351] = 24'b000010011000011011011001;
        rom[1352] = 24'b000011010111000000111000;
        rom[1353] = 24'b000011101000010010111001;
        rom[1354] = 24'b000010110101011111110100;
        rom[1355] = 24'b000001111011010101111011;
        rom[1356] = 24'b000001111101010111010101;
        rom[1357] = 24'b000010110111100010101100;
        rom[1358] = 24'b000011110000011101011011;
        rom[1359] = 24'b000011011010111100001000;
        rom[1360] = 24'b000010010110000001011110;
        rom[1361] = 24'b000001110010111110100111;
        rom[1362] = 24'b000010001110110100101000;
        rom[1363] = 24'b000011011010000111010010;
        rom[1364] = 24'b000011110000110001011001;
        rom[1365] = 24'b000011000010000001010000;
        rom[1366] = 24'b000010000101111010001000;
        rom[1367] = 24'b000010000100101010111111;
        rom[1368] = 24'b000010111110011011100000;
        rom[1369] = 24'b000011110000110111010000;
        rom[1370] = 24'b000011100101110111000111;
        rom[1371] = 24'b000010100010011011001111;
        rom[1372] = 24'b000001101100010110010110;
        rom[1373] = 24'b000010001111001101101101;
        rom[1374] = 24'b000011010011001011101000;
        rom[1375] = 24'b000011110001011101111000;
        rom[1376] = 24'b000011000010001101110001;
        rom[1377] = 24'b000001111101010011000111;
        rom[1378] = 24'b000001101010001110000100;
        rom[1379] = 24'b000010100011001000110011;
        rom[1380] = 24'b000011100010001100101010;
        rom[1381] = 24'b000011011100111001010100;
        rom[1382] = 24'b000010011000111110011011;
        rom[1383] = 24'b000001101011000011110110;
        rom[1384] = 24'b000001111001111001100111;
        rom[1385] = 24'b000011000010010000000110;
        rom[1386] = 24'b000011100101011111100000;
        rom[1387] = 24'b000011000100101100010110;
        rom[1388] = 24'b000010000110000110110111;
        rom[1389] = 24'b000001101000100111100110;
        rom[1390] = 24'b000010011000111110011011;
        rom[1391] = 24'b000011010000101100000100;
        rom[1392] = 24'b000011011000011011101010;
        rom[1393] = 24'b000010100011001000110011;
        rom[1394] = 24'b000001101100101010010100;
        rom[1395] = 24'b000010000010001011100111;
        rom[1396] = 24'b000010111000011100110001;
        rom[1397] = 24'b000011100010110100011000;
        rom[1398] = 24'b000011000100100010000111;
        rom[1399] = 24'b000010000011000000011101;
        rom[1400] = 24'b000001101001111010000110;
        rom[1401] = 24'b000010010011110001101111;
        rom[1402] = 24'b000011001111111000110111;
        rom[1403] = 24'b000011011101010101010000;
        rom[1404] = 24'b000010101010111001011111;
        rom[1405] = 24'b000001110110000001011111;
        rom[1406] = 24'b000001111001101100111000;
        rom[1407] = 24'b000010110011010111110000;
        rom[1408] = 24'b000011010101111010101001;
        rom[1409] = 24'b000011000001101100110010;
        rom[1410] = 24'b000010000010100111010111;
        rom[1411] = 24'b000001100110110001010111;
        rom[1412] = 24'b000010010110000001011110;
        rom[1413] = 24'b000011010011100111011000;
        rom[1414] = 24'b000011010101100110101011;
        rom[1415] = 24'b000010101011010101011100;
        rom[1416] = 24'b000001111000011110110101;
        rom[1417] = 24'b000001111011010101111011;
        rom[1418] = 24'b000010110000100111010100;
        rom[1419] = 24'b000011100000111110001001;
        rom[1420] = 24'b000011001010110011101000;
        rom[1421] = 24'b000010001001110001111001;
        rom[1422] = 24'b000001101000111110110000;
        rom[1423] = 24'b000010001100001110001001;
        rom[1424] = 24'b000011001101001111111000;
        rom[1425] = 24'b000011011100000101101001;
        rom[1426] = 24'b000010101011101110110100;
        rom[1427] = 24'b000001101111001000101011;
        rom[1428] = 24'b000001110011100110010101;
        rom[1429] = 24'b000010101101110001101100;
        rom[1430] = 24'b000011100001110011111011;
        rom[1431] = 24'b000011001001110110011000;
        rom[1432] = 24'b000010000111010111111110;
        rom[1433] = 24'b000001100100010101000111;
        rom[1434] = 24'b000010000111011111111000;
        rom[1435] = 24'b000011001101111010000010;
        rom[1436] = 24'b000011101011111000111001;
        rom[1437] = 24'b000011000010000001010000;
        rom[1438] = 24'b000010000011011101111000;
        rom[1439] = 24'b000010001001100011011111;
        rom[1440] = 24'b000011000011010100000000;
        rom[1441] = 24'b000100000001111101000000;
        rom[1442] = 24'b000011110110111100110111;
        rom[1443] = 24'b000010110101111101001111;
        rom[1444] = 24'b000010001100000101100110;
        rom[1445] = 24'b000010101010000100011101;
        rom[1446] = 24'b000011110010111010110111;
        rom[1447] = 24'b000100010001001101001000;
        rom[1448] = 24'b000011110000100110100001;
        rom[1449] = 24'b000010101001001111100111;
        rom[1450] = 24'b000010011011000011000100;
        rom[1451] = 24'b000011010110011010000011;
        rom[1452] = 24'b000100001011101100111010;
        rom[1453] = 24'b000100001011010010000100;
        rom[1454] = 24'b000011001001110011011011;
        rom[1455] = 24'b000010010100100100000110;
        rom[1456] = 24'b000010100011011001110111;
        rom[1457] = 24'b000011101011110000010110;
        rom[1458] = 24'b000100010011111000010000;
        rom[1459] = 24'b000011110000101000110110;
        rom[1460] = 24'b000010100101110110000111;
        rom[1461] = 24'b000010001111101011100110;
        rom[1462] = 24'b000011000010011110101011;
        rom[1463] = 24'b000100001000110101110100;
        rom[1464] = 24'b000100010111111010001010;
        rom[1465] = 24'b000011100010100111010011;
        rom[1466] = 24'b000010100111010000010100;
        rom[1467] = 24'b000010101011101011110111;
        rom[1468] = 24'b000011011000001100000001;
        rom[1469] = 24'b000100000000000111011000;
        rom[1470] = 24'b000011011010100000010111;
        rom[1471] = 24'b000010011000111110101101;
        rom[1472] = 24'b000001110011101011000110;
        rom[1473] = 24'b000010010110001101111111;
        rom[1474] = 24'b000011001111111000110111;
        rom[1475] = 24'b000011011000011100110000;
        rom[1476] = 24'b000010011110101100001111;
        rom[1477] = 24'b000001100100111011101111;
        rom[1478] = 24'b000001101101011111101000;
        rom[1479] = 24'b000010110000111011100000;
        rom[1480] = 24'b000011010101111010101001;
        rom[1481] = 24'b000011000001101100110010;
        rom[1482] = 24'b000010000010100111010111;
        rom[1483] = 24'b000001100100010101000111;
        rom[1484] = 24'b000010001001110100001110;
        rom[1485] = 24'b000011000100111101111000;
        rom[1486] = 24'b000011001011110101101011;
        rom[1487] = 24'b000010011111001000001100;
        rom[1488] = 24'b000001011101101000000101;
        rom[1489] = 24'b000001101100101100011011;
        rom[1490] = 24'b000010101011101110110100;
        rom[1491] = 24'b000011010010010100101001;
        rom[1492] = 24'b000010110100110101011000;
        rom[1493] = 24'b000001111101100100101001;
        rom[1494] = 24'b000001100001101010000000;
        rom[1495] = 24'b000010000010011101001001;
        rom[1496] = 24'b000011000011011110111000;
        rom[1497] = 24'b000011010100110000111001;
        rom[1498] = 24'b000010011000001100110100;
        rom[1499] = 24'b000001010110101110001011;
        rom[1500] = 24'b000001010001011010110101;
        rom[1501] = 24'b000001111100111100101100;
        rom[1502] = 24'b000010100010010101011011;
        rom[1503] = 24'b000010001010010111111000;
        rom[1504] = 24'b000000111001001111111110;
        rom[1505] = 24'b000000000000001110110111;
        rom[1506] = 24'b000000100000111101010111;
        rom[1507] = 24'b000001111000011101010010;
        rom[1508] = 24'b000010111101100000001001;
        rom[1509] = 24'b000011000110111001110000;
        rom[1510] = 24'b000011001010010001001000;
        rom[1511] = 24'b000100100011010111001111;
        rom[1512] = 24'b000111100000111101010000;
        rom[1513] = 24'b001010100000111111100000;
        rom[1514] = 24'b001011111100100001110111;
        rom[1515] = 24'b001011100111011110101111;
        rom[1516] = 24'b001010001111001110010110;
        rom[1517] = 24'b001000100010000010111101;
        rom[1518] = 24'b000110100101001001001000;
        rom[1519] = 24'b000100011010111110001000;
        rom[1520] = 24'b000010001100100000010001;
        rom[1521] = 24'b000000100111110110010111;
        rom[1522] = 24'b000000011110100010010100;
        rom[1523] = 24'b000001100110000110100011;
        rom[1524] = 24'b000010111000101100011010;
        rom[1525] = 24'b000010111010101101110100;
        rom[1526] = 24'b000001111011101011011011;
        rom[1527] = 24'b000001001011010100100110;
        rom[1528] = 24'b000001011100100110100111;
        rom[1529] = 24'b000010100010100000110110;
        rom[1530] = 24'b000011001010101000110000;
        rom[1531] = 24'b000010100100111101000110;
        rom[1532] = 24'b000001100011111011010111;
        rom[1533] = 24'b000001001000111000010110;
        rom[1534] = 24'b000001110100010110101011;
        rom[1535] = 24'b000010110000111100110100;
        rom[1536] = 24'b000010111101100100111010;
        rom[1537] = 24'b000010000011011001100011;
        rom[1538] = 24'b000001001000000010100100;
        rom[1539] = 24'b000001010110001111000111;
        rom[1540] = 24'b000010010001011000110001;
        rom[1541] = 24'b000010111011110000011000;
        rom[1542] = 24'b000010100100110010110111;
        rom[1543] = 24'b000001100011010001001101;
        rom[1544] = 24'b000001000111101110100110;
        rom[1545] = 24'b000001101100101101101111;
        rom[1546] = 24'b000010101011010001000111;
        rom[1547] = 24'b000010110011110101000000;
        rom[1548] = 24'b000010000011110101100000;
        rom[1549] = 24'b000001010001011001101111;
        rom[1550] = 24'b000001011001111101101000;
        rom[1551] = 24'b000010001110110000000000;
        rom[1552] = 24'b000010111000100111101001;
        rom[1553] = 24'b000010100100011001110010;
        rom[1554] = 24'b000001100111110000100111;
        rom[1555] = 24'b000001001001011110010111;
        rom[1556] = 24'b000001110001011001101110;
        rom[1557] = 24'b000010101100100011011000;
        rom[1558] = 24'b000010111000010011101011;
        rom[1559] = 24'b000010000100010001011100;
        rom[1560] = 24'b000001001110111110100101;
        rom[1561] = 24'b000001010110101110001011;
        rom[1562] = 24'b000010010000111000000100;
        rom[1563] = 24'b000010111001111010001001;
        rom[1564] = 24'b000010011110110111001000;
        rom[1565] = 24'b000001100010101101111001;
        rom[1566] = 24'b000001000100010111000000;
        rom[1567] = 24'b000001100101001010001001;
        rom[1568] = 24'b000010101000101000001000;
        rom[1569] = 24'b000010110111011101111001;
        rom[1570] = 24'b000010000010001110100100;
        rom[1571] = 24'b000001000101101000011011;
        rom[1572] = 24'b000001001010000110000101;
        rom[1573] = 24'b000010001011100110001100;
        rom[1574] = 24'b000011000010000100101011;
        rom[1575] = 24'b000010101110111111101000;
        rom[1576] = 24'b000001101010000100111110;
        rom[1577] = 24'b000001000010001001100111;
        rom[1578] = 24'b000001100101010100011000;
        rom[1579] = 24'b000010101011101110100010;
        rom[1580] = 24'b000010111011000011111001;
        rom[1581] = 24'b000010001001110111100000;
        rom[1582] = 24'b000001001011010100001000;
        rom[1583] = 24'b000001000101001100011111;
        rom[1584] = 24'b000001111100100000110000;
        rom[1585] = 24'b000010111000101101100000;
        rom[1586] = 24'b000010101000110100110111;
        rom[1587] = 24'b000001101100101101101111;
        rom[1588] = 24'b000000111011100001010110;
        rom[1589] = 24'b000001011011111100011101;
        rom[1590] = 24'b000010100010010110101000;
        rom[1591] = 24'b000010111110001100101000;
        rom[1592] = 24'b000010011000101101100001;
        rom[1593] = 24'b000001011000101011010111;
        rom[1594] = 24'b000001000101100110010100;
        rom[1595] = 24'b000001111110100001000011;
        rom[1596] = 24'b000010111011001000101010;
        rom[1597] = 24'b000010111000010001100100;
        rom[1598] = 24'b000001110110110010111011;
        rom[1599] = 24'b000001000011111111110110;
        rom[1600] = 24'b000001010000011001010111;
        rom[1601] = 24'b000010010001011011000110;
        rom[1602] = 24'b000010111011111111010000;
        rom[1603] = 24'b000010011000101111110110;
        rom[1604] = 24'b000001010010110101100111;
        rom[1605] = 24'b000000111010001110110110;
        rom[1606] = 24'b000001100011010000111011;
        rom[1607] = 24'b000010100010010011010100;
        rom[1608] = 24'b000010100111100110101010;
        rom[1609] = 24'b000001101111110111100011;
        rom[1610] = 24'b000000111011110101010100;
        rom[1611] = 24'b000001000000010000110111;
        rom[1612] = 24'b000010000010101111010001;
        rom[1613] = 24'b000010101010101010101000;
        rom[1614] = 24'b000010010001010000110111;
        rom[1615] = 24'b000001001111101111001101;
        rom[1616] = 24'b000000110001110000010110;
        rom[1617] = 24'b000001100000100000011111;
        rom[1618] = 24'b000010011010001011010111;
        rom[1619] = 24'b000010101100100000010000;
        rom[1620] = 24'b000001110101001011111111;
        rom[1621] = 24'b000001000101001100011111;
        rom[1622] = 24'b000001010101000101001000;
        rom[1623] = 24'b000010010011101000100000;
        rom[1624] = 24'b000011000111010001001001;
        rom[1625] = 24'b000010110111111011110010;
        rom[1626] = 24'b000010000101000011100111;
        rom[1627] = 24'b000001101001001101100111;
        rom[1628] = 24'b000010010011100101001110;
        rom[1629] = 24'b000011010001001011001000;
        rom[1630] = 24'b000011011111010111101011;
        rom[1631] = 24'b000010110101000110011100;
        rom[1632] = 24'b000010000010001111110101;
        rom[1633] = 24'b000010001001111111011011;
        rom[1634] = 24'b000011000100001001010100;
        rom[1635] = 24'b000011110100100000001001;
        rom[1636] = 24'b000011010111000000111000;
        rom[1637] = 24'b000010011101010011111001;
        rom[1638] = 24'b000001111110111101000000;
        rom[1639] = 24'b000010100100101000101001;
        rom[1640] = 24'b000011011011111001011000;
        rom[1641] = 24'b000011110100100000001001;
        rom[1642] = 24'b000011000001101101000100;
        rom[1643] = 24'b000010000111100011001011;
        rom[1644] = 24'b000010001001100100100101;
        rom[1645] = 24'b000011000110001100001100;
        rom[1646] = 24'b000011111010001110011011;
        rom[1647] = 24'b000011100100101101001000;
        rom[1648] = 24'b000010100100101010111110;
        rom[1649] = 24'b000001111111001011110111;
        rom[1650] = 24'b000010100100110010111000;
        rom[1651] = 24'b000011100110010100100010;
        rom[1652] = 24'b000011111111011010111001;
        rom[1653] = 24'b000011010000101010110000;
        rom[1654] = 24'b000010001010110010101000;
        rom[1655] = 24'b000010000100101010111111;
        rom[1656] = 24'b000011000000110111101111;
        rom[1657] = 24'b000011111000001100000000;
        rom[1658] = 24'b000011101000010011010111;
        rom[1659] = 24'b000010100111010011101111;
        rom[1660] = 24'b000001110110000111010110;
        rom[1661] = 24'b000010010100000110001101;
        rom[1662] = 24'b000011010101100111111000;
        rom[1663] = 24'b000011111000110010101000;
        rom[1664] = 24'b000011001110011011000001;
        rom[1665] = 24'b000010001001100000010111;
        rom[1666] = 24'b000001111000110111100100;
        rom[1667] = 24'b000010101010011101100011;
        rom[1668] = 24'b000011101011111101101010;
        rom[1669] = 24'b000011100110101010010100;
        rom[1670] = 24'b000010100111100111111011;
        rom[1671] = 24'b000001110100110100110110;
        rom[1672] = 24'b000010000001001110010111;
        rom[1673] = 24'b000011000010010000000110;
        rom[1674] = 24'b000011101010011000000000;
        rom[1675] = 24'b000011001001100100110110;
        rom[1676] = 24'b000010000110000110110111;
        rom[1677] = 24'b000001110010011000100110;
        rom[1678] = 24'b000010011101110110111011;
        rom[1679] = 24'b000011011100111001010100;
        rom[1680] = 24'b000011100100101000111010;
        rom[1681] = 24'b000010100101100101000011;
        rom[1682] = 24'b000001110011111111000100;
        rom[1683] = 24'b000001111010110110110111;
        rom[1684] = 24'b000010111010111001000001;
        rom[1685] = 24'b000011100111101100111000;
        rom[1686] = 24'b000011001110010011000111;
        rom[1687] = 24'b000010001100110001011101;
        rom[1688] = 24'b000001110011101011000110;
        rom[1689] = 24'b000010010110001101111111;
        rom[1690] = 24'b000011010010010101000111;
        rom[1691] = 24'b000011011101010101010000;
        rom[1692] = 24'b000010101010111001011111;
        rom[1693] = 24'b000001110001001000111111;
        rom[1694] = 24'b000001111001101100111000;
        rom[1695] = 24'b000010110101110100000000;
        rom[1696] = 24'b000011011111101011101001;
        rom[1697] = 24'b000011001001000001100010;
        rom[1698] = 24'b000010001001111100000111;
        rom[1699] = 24'b000001101011101001110111;
        rom[1700] = 24'b000010010110000001011110;
        rom[1701] = 24'b000011010011100111011000;
        rom[1702] = 24'b000011011111010111101011;
        rom[1703] = 24'b000010101101110001101100;
        rom[1704] = 24'b000001111000011110110101;
        rom[1705] = 24'b000010000000001110011011;
        rom[1706] = 24'b000010110011000011100100;
        rom[1707] = 24'b000011101000010010111001;
        rom[1708] = 24'b000011001010110011101000;
        rom[1709] = 24'b000010001100001110001001;
        rom[1710] = 24'b000001110010101111110000;
        rom[1711] = 24'b000010010001000110101001;
        rom[1712] = 24'b000011001101001111111000;
        rom[1713] = 24'b000011100000111110001001;
        rom[1714] = 24'b000010101110001011000100;
        rom[1715] = 24'b000001110100000001001011;
        rom[1716] = 24'b000001110001001010000101;
        rom[1717] = 24'b000010110000001101111100;
        rom[1718] = 24'b000011100100010000001011;
        rom[1719] = 24'b000011010001001011001000;
        rom[1720] = 24'b000010010001001000111110;
        rom[1721] = 24'b000001101011101001110111;
        rom[1722] = 24'b000010001110110100101000;
        rom[1723] = 24'b000011010000010110010010;
        rom[1724] = 24'b000011101001011100101001;
        rom[1725] = 24'b000010110101110100000000;
        rom[1726] = 24'b000001110111010000101000;
        rom[1727] = 24'b000001110011100101001111;
        rom[1728] = 24'b000010101101010101110000;
        rom[1729] = 24'b000011101001100010100000;
        rom[1730] = 24'b000011100000111110100111;
        rom[1731] = 24'b000010100111010011101111;
        rom[1732] = 24'b000001110001001110110110;
        rom[1733] = 24'b000010010001101001111101;
        rom[1734] = 24'b000011011111011000111000;
        rom[1735] = 24'b000100000111011100001000;
        rom[1736] = 24'b000011011111100000110001;
        rom[1737] = 24'b000010011101000010010111;
        rom[1738] = 24'b000010001100011001100100;
        rom[1739] = 24'b000011000101010100010011;
        rom[1740] = 24'b000100001001010000101010;
        rom[1741] = 24'b000100001000110101110100;
        rom[1742] = 24'b000011001110101011111011;
        rom[1743] = 24'b000010100000110001010110;
        rom[1744] = 24'b000010110100011111100111;
        rom[1745] = 24'b000011110111111101100110;
        rom[1746] = 24'b000100100010100001110000;
        rom[1747] = 24'b000011111100110110000110;
        rom[1748] = 24'b000010111011110100010111;
        rom[1749] = 24'b000010011110010101000110;
        rom[1750] = 24'b000011001001110011011011;
        rom[1751] = 24'b000100000011111101010100;
        rom[1752] = 24'b000100001011101100111010;
        rom[1753] = 24'b000011011000110110010011;
        rom[1754] = 24'b000010011000100110110100;
        rom[1755] = 24'b000010100110110011010111;
        rom[1756] = 24'b000011100001111101000001;
        rom[1757] = 24'b000100010001001101001000;
        rom[1758] = 24'b000011111111001000001000;
        rom[1759] = 24'b000011000010011110111101;
        rom[1760] = 24'b000010011111100111100110;
        rom[1761] = 24'b000010111010110101101111;
        rom[1762] = 24'b000011101111101000000111;
        rom[1763] = 24'b000011110011010011100000;
        rom[1764] = 24'b000010110100101010011111;
        rom[1765] = 24'b000001111010111001111111;
        rom[1766] = 24'b000001111100001001001000;
        rom[1767] = 24'b000010110101110100000000;
        rom[1768] = 24'b000011100100100100001001;
        rom[1769] = 24'b000011001101111010000010;
        rom[1770] = 24'b000010000111011111110111;
        rom[1771] = 24'b000001101001001101100111;
        rom[1772] = 24'b000010001110101100101110;
        rom[1773] = 24'b000011001100010010101000;
        rom[1774] = 24'b000011011000000010111011;
        rom[1775] = 24'b000010100110011100111100;
        rom[1776] = 24'b000001101110101101110101;
        rom[1777] = 24'b000001111000111001101011;
        rom[1778] = 24'b000010110011000011100100;
        rom[1779] = 24'b000011011110100001111001;
        rom[1780] = 24'b000011000101111011001000;
        rom[1781] = 24'b000010000100111001011001;
        rom[1782] = 24'b000001100001101010000000;
        rom[1783] = 24'b000010001001110001111001;
        rom[1784] = 24'b000011001000010111011000;
        rom[1785] = 24'b000011011001101001011001;
        rom[1786] = 24'b000010100100011010000100;
        rom[1787] = 24'b000001101111001000101011;
        rom[1788] = 24'b000001101100010001100101;
        rom[1789] = 24'b000010100110011100111100;
        rom[1790] = 24'b000011011010011111001011;
        rom[1791] = 24'b000011001001110110011000;
        rom[1792] = 24'b000010000100111011101110;
        rom[1793] = 24'b000001011000000111110111;
        rom[1794] = 24'b000001110011111101111000;
        rom[1795] = 24'b000010100100011001110010;
        rom[1796] = 24'b000010101001111110001001;
        rom[1797] = 24'b000001101100100100100000;
        rom[1798] = 24'b000000100110101100011000;
        rom[1799] = 24'b000000010001111011001111;
        rom[1800] = 24'b000001000001111010101111;
        rom[1801] = 24'b000010000111111000100000;
        rom[1802] = 24'b000010101011010001000111;
        rom[1803] = 24'b000010101110101000011111;
        rom[1804] = 24'b000011001001000111110110;
        rom[1805] = 24'b000101000011111000001101;
        rom[1806] = 24'b000111111000001001100111;
        rom[1807] = 24'b001010011111001001111000;
        rom[1808] = 24'b001011100111100010000001;
        rom[1809] = 24'b001011101001011010100111;
        rom[1810] = 24'b001011001111000000110100;
        rom[1811] = 24'b001010111100001111110011;
        rom[1812] = 24'b001001010101010010101010;
        rom[1813] = 24'b000110000010111010010100;
        rom[1814] = 24'b000010101100100000011011;
        rom[1815] = 24'b000000110010111010000110;
        rom[1816] = 24'b000000111010011011000111;
        rom[1817] = 24'b000010010001011011000110;
        rom[1818] = 24'b000011001010101000110000;
        rom[1819] = 24'b000010110001001010010110;
        rom[1820] = 24'b000001110000001000100111;
        rom[1821] = 24'b000001010111100001110110;
        rom[1822] = 24'b000010000011000000001011;
        rom[1823] = 24'b000010111111100110010100;
        rom[1824] = 24'b000011000100111001101010;
        rom[1825] = 24'b000010001101001010100011;
        rom[1826] = 24'b000001011011100100100100;
        rom[1827] = 24'b000001100111010100110111;
        rom[1828] = 24'b000010100000000010010001;
        rom[1829] = 24'b000011000111111101101000;
        rom[1830] = 24'b000010101110100011111000;
        rom[1831] = 24'b000001101111011110011101;
        rom[1832] = 24'b000001010110011000000110;
        rom[1833] = 24'b000001111011010111001111;
        rom[1834] = 24'b000010110101000010000111;
        rom[1835] = 24'b000011000010011110100000;
        rom[1836] = 24'b000010001011001010010000;
        rom[1837] = 24'b000001010001011001101111;
        rom[1838] = 24'b000001011100011001111000;
        rom[1839] = 24'b000010010110000100110000;
        rom[1840] = 24'b000010111011000011111001;
        rom[1841] = 24'b000010100110110110000010;
        rom[1842] = 24'b000001100111110000101000;
        rom[1843] = 24'b000001010000110011000111;
        rom[1844] = 24'b000001110001011001101110;
        rom[1845] = 24'b000010110001011011111000;
        rom[1846] = 24'b000010111101001100001011;
        rom[1847] = 24'b000010001001001001111100;
        rom[1848] = 24'b000001010001011010110101;
        rom[1849] = 24'b000001010110101110001011;
        rom[1850] = 24'b000010010011010100010100;
        rom[1851] = 24'b000011000001001110111001;
        rom[1852] = 24'b000010101000101000001000;
        rom[1853] = 24'b000001101110111011001001;
        rom[1854] = 24'b000001001110001000000000;
        rom[1855] = 24'b000001110110001111111001;
        rom[1856] = 24'b000010110111010001101000;
        rom[1857] = 24'b000011001000100011101001;
        rom[1858] = 24'b000010010011010100010100;
        rom[1859] = 24'b000001011001001010011011;
        rom[1860] = 24'b000001011101101000000101;
        rom[1861] = 24'b000010010111110011011100;
        rom[1862] = 24'b000011001011110101101011;
        rom[1863] = 24'b000010111011001100111000;
        rom[1864] = 24'b000001110110010010001110;
        rom[1865] = 24'b000001010101101011100111;
        rom[1866] = 24'b000001101010001100110111;
        rom[1867] = 24'b000010110011000011010010;
        rom[1868] = 24'b000011001110100101111001;
        rom[1869] = 24'b000010011101011001100000;
        rom[1870] = 24'b000001011001111101101000;
        rom[1871] = 24'b000001010001011001101111;
        rom[1872] = 24'b000010001011001010001111;
        rom[1873] = 24'b000011000111010111000000;
        rom[1874] = 24'b000010111110110011000111;
        rom[1875] = 24'b000001111011010111001111;
        rom[1876] = 24'b000001001010001010110110;
        rom[1877] = 24'b000001100101101101011101;
        rom[1878] = 24'b000010101001101011010111;
        rom[1879] = 24'b000011001100110110001000;
        rom[1880] = 24'b000010100010011110100001;
        rom[1881] = 24'b000001100000000000000111;
        rom[1882] = 24'b000001001111010111010100;
        rom[1883] = 24'b000010001000010010000011;
        rom[1884] = 24'b000011000010011101011010;
        rom[1885] = 24'b000011000100011110110100;
        rom[1886] = 24'b000010000111111000101011;
        rom[1887] = 24'b000001011001111110000110;
        rom[1888] = 24'b000001100001011111000111;
        rom[1889] = 24'b000010101110101110000110;
        rom[1890] = 24'b000011010001111101100000;
        rom[1891] = 24'b000010110001001010010110;
        rom[1892] = 24'b000001101000110011110111;
        rom[1893] = 24'b000001010010101001010110;
        rom[1894] = 24'b000001111001001111001011;
        rom[1895] = 24'b000010111010101101110100;
        rom[1896] = 24'b000011000100111001101010;
        rom[1897] = 24'b000010001010101110010011;
        rom[1898] = 24'b000001011001001000010100;
        rom[1899] = 24'b000001100000000000000111;
        rom[1900] = 24'b000010011101100110000001;
        rom[1901] = 24'b000011000101100001011000;
        rom[1902] = 24'b000010100111001111001000;
        rom[1903] = 24'b000001100101101101011101;
        rom[1904] = 24'b000001010011111011110110;
        rom[1905] = 24'b000001111011010111001111;
        rom[1906] = 24'b000010110101000010000111;
        rom[1907] = 24'b000011000100111010110000;
        rom[1908] = 24'b000010010010011111000000;
        rom[1909] = 24'b000001011000101110011111;
        rom[1910] = 24'b000001100001010010011000;
        rom[1911] = 24'b000010011000100001000000;
        rom[1912] = 24'b000010111101100000001001;
        rom[1913] = 24'b000010110011000011010010;
        rom[1914] = 24'b000001110011111101111000;
        rom[1915] = 24'b000001011010100100000111;
        rom[1916] = 24'b000001111011001010101110;
        rom[1917] = 24'b000010110110010100011000;
        rom[1918] = 24'b000011000110111101001011;
        rom[1919] = 24'b000010010111110011011100;
        rom[1920] = 24'b000001100010100000100101;
        rom[1921] = 24'b000001101100101100011011;
        rom[1922] = 24'b000010101001010010100100;
        rom[1923] = 24'b000011100000111110001001;
        rom[1924] = 24'b000011001101001111111000;
        rom[1925] = 24'b000010010011100010111001;
        rom[1926] = 24'b000001110010101111110000;
        rom[1927] = 24'b000010011101010011111001;
        rom[1928] = 24'b000011100011001110001000;
        rom[1929] = 24'b000011110110111100011001;
        rom[1930] = 24'b000011000001101101000100;
        rom[1931] = 24'b000010001100011011101011;
        rom[1932] = 24'b000010001110011101000101;
        rom[1933] = 24'b000011000011101111111100;
        rom[1934] = 24'b000011110111110010001011;
        rom[1935] = 24'b000011101001100101101000;
        rom[1936] = 24'b000010100100101010111110;
        rom[1937] = 24'b000001111100101111100111;
        rom[1938] = 24'b000010011111111010010111;
        rom[1939] = 24'b000011100011111000010010;
        rom[1940] = 24'b000011111010100010011001;
        rom[1941] = 24'b000011001011110010010000;
        rom[1942] = 24'b000010001010110010101000;
        rom[1943] = 24'b000010000010001110101111;
        rom[1944] = 24'b000010111110011011011111;
        rom[1945] = 24'b000011110101101111110000;
        rom[1946] = 24'b000011101010101111100111;
        rom[1947] = 24'b000010101001101111111111;
        rom[1948] = 24'b000001111000100011100110;
        rom[1949] = 24'b000010010100000110001101;
        rom[1950] = 24'b000011011010100000010111;
        rom[1951] = 24'b000011111011001110111000;
        rom[1952] = 24'b000011010000110111010001;
        rom[1953] = 24'b000010010000110101000111;
        rom[1954] = 24'b000001111101110000000100;
        rom[1955] = 24'b000010110110101010110011;
        rom[1956] = 24'b000011110011010010011010;
        rom[1957] = 24'b000011110010110111100100;
        rom[1958] = 24'b000010110011110101001011;
        rom[1959] = 24'b000001111110100101110110;
        rom[1960] = 24'b000010001000100011000111;
        rom[1961] = 24'b000011001100000001000110;
        rom[1962] = 24'b000011111001000001100000;
        rom[1963] = 24'b000011011101000110110110;
        rom[1964] = 24'b000010011100000101000111;
        rom[1965] = 24'b000010000101111010100110;
        rom[1966] = 24'b000010110001011000111011;
        rom[1967] = 24'b000011101101111111000100;
        rom[1968] = 24'b000011111000001010111010;
        rom[1969] = 24'b000011000000011011110011;
        rom[1970] = 24'b000010001100011001100100;
        rom[1971] = 24'b000010011010100110000111;
        rom[1972] = 24'b000011010011010011100001;
        rom[1973] = 24'b000100000010100011101000;
        rom[1974] = 24'b000011101110000010011000;
        rom[1975] = 24'b000010110001011001001101;
        rom[1976] = 24'b000010011000010010110110;
        rom[1977] = 24'b000010111101010001111111;
        rom[1978] = 24'b000011111011110101010111;
        rom[1979] = 24'b000100000110110101100000;
        rom[1980] = 24'b000011011110001010110000;
        rom[1981] = 24'b000010100100011010001111;
        rom[1982] = 24'b000010100000110000111000;
        rom[1983] = 24'b000011011010011011110000;
        rom[1984] = 24'b000100010010111100111001;
        rom[1985] = 24'b000100000110000011110010;
        rom[1986] = 24'b000011000010000101111000;
        rom[1987] = 24'b000010011110111011000111;
        rom[1988] = 24'b000011000001111101111110;
        rom[1989] = 24'b000011111101000111101000;
        rom[1990] = 24'b000100001011010100001011;
        rom[1991] = 24'b000011010100110101101100;
        rom[1992] = 24'b000010011000001110000101;
        rom[1993] = 24'b000010010001010100001011;
        rom[1994] = 24'b000011000110100101100100;
        rom[1995] = 24'b000011101000010010111001;
        rom[1996] = 24'b000011010010001000011000;
        rom[1997] = 24'b000010010001000110101001;
        rom[1998] = 24'b000001110010101111110000;
        rom[1999] = 24'b000010001100001110001001;
        rom[2000] = 24'b000011001000010111011000;
        rom[2001] = 24'b000011011001101001011001;
        rom[2002] = 24'b000010100001111101110100;
        rom[2003] = 24'b000001100010111011011011;
        rom[2004] = 24'b000001100010100000100101;
        rom[2005] = 24'b000010100001100100011100;
        rom[2006] = 24'b000011010011001010011011;
        rom[2007] = 24'b000010111011001100111000;
        rom[2008] = 24'b000001110110010010001110;
        rom[2009] = 24'b000001010011001111010111;
        rom[2010] = 24'b000001110011111101110111;
        rom[2011] = 24'b000010110111111011110010;
        rom[2012] = 24'b000011010001000010001001;
        rom[2013] = 24'b000010100010010010000000;
        rom[2014] = 24'b000001011110110110001000;
        rom[2015] = 24'b000001100000000011001111;
        rom[2016] = 24'b000010011100001111111111;
        rom[2017] = 24'b000011010001001000000000;
        rom[2018] = 24'b000011001000100100000111;
        rom[2019] = 24'b000010001100011100111111;
        rom[2020] = 24'b000001011000110100010110;
        rom[2021] = 24'b000001111001001111011101;
        rom[2022] = 24'b000010111010110001000111;
        rom[2023] = 24'b000011011101111011111000;
        rom[2024] = 24'b000010101110101011110001;
        rom[2025] = 24'b000001110001000101110111;
        rom[2026] = 24'b000001010110101100000100;
        rom[2027] = 24'b000010001111100110110011;
        rom[2028] = 24'b000011000100111001101010;
        rom[2029] = 24'b000010110101110101010100;
        rom[2030] = 24'b000001101010100101101011;
        rom[2031] = 24'b000000100100010000100110;
        rom[2032] = 24'b000000100010000000100111;
        rom[2033] = 24'b000001100011000010010110;
        rom[2034] = 24'b000001110111101000010000;
        rom[2035] = 24'b000001001010100111110110;
        rom[2036] = 24'b000000011000001111100111;
        rom[2037] = 24'b000000110010111010000110;
        rom[2038] = 24'b000010100111100111111011;
        rom[2039] = 24'b000100110100110010010100;
        rom[2040] = 24'b000110001000001101101010;
        rom[2041] = 24'b000111000000110010000011;
        rom[2042] = 24'b001000000110110100010100;
        rom[2043] = 24'b001010000010111000000111;
        rom[2044] = 24'b001011111000100111110001;
        rom[2045] = 24'b001100101111001100101000;
        rom[2046] = 24'b001011001100100011011000;
        rom[2047] = 24'b000111100111011100111101;
        rom[2048] = 24'b000011111110110101010110;
        rom[2049] = 24'b000010010011110001101111;
        rom[2050] = 24'b000010001011100001110111;
        rom[2051] = 24'b000010011000111110010000;
        rom[2052] = 24'b000001111100100000110000;
        rom[2053] = 24'b000001011000101110011111;
        rom[2054] = 24'b000001100110001010111000;
        rom[2055] = 24'b000010011010111101010000;
        rom[2056] = 24'b000010111111111100011001;
        rom[2057] = 24'b000010110000100111000010;
        rom[2058] = 24'b000001101010001100111000;
        rom[2059] = 24'b000001010011001111010111;
        rom[2060] = 24'b000001110110010010001110;
        rom[2061] = 24'b000010110001011011111000;
        rom[2062] = 24'b000010111010101111111011;
        rom[2063] = 24'b000010001110000010011100;
        rom[2064] = 24'b000001011000101111100101;
        rom[2065] = 24'b000001011001001010011011;
        rom[2066] = 24'b000010010101110000100100;
        rom[2067] = 24'b000011000001001110111001;
        rom[2068] = 24'b000010101011000100011000;
        rom[2069] = 24'b000001100111100110011001;
        rom[2070] = 24'b000001000110110011010000;
        rom[2071] = 24'b000001101110111011001001;
        rom[2072] = 24'b000010101111111100111000;
        rom[2073] = 24'b000011000001001110111001;
        rom[2074] = 24'b000010001110011011110100;
        rom[2075] = 24'b000001010110101110001011;
        rom[2076] = 24'b000001010110010011010101;
        rom[2077] = 24'b000010001110000010011100;
        rom[2078] = 24'b000011000100100000111011;
        rom[2079] = 24'b000010101010000111001000;
        rom[2080] = 24'b000001100101001100011110;
        rom[2081] = 24'b000001000100100101110111;
        rom[2082] = 24'b000001100000011011110111;
        rom[2083] = 24'b000010101011101110100010;
        rom[2084] = 24'b000011000100110100111001;
        rom[2085] = 24'b000010011000100001000000;
        rom[2086] = 24'b000001010101000101001000;
        rom[2087] = 24'b000001001100100001001111;
        rom[2088] = 24'b000010001000101101111111;
        rom[2089] = 24'b000011000111010111000000;
        rom[2090] = 24'b000010111100010110110111;
        rom[2091] = 24'b000001110110011110101111;
        rom[2092] = 24'b000001000111101110100110;
        rom[2093] = 24'b000001100101101101011101;
        rom[2094] = 24'b000010100010010110100111;
        rom[2095] = 24'b000011000101100001011000;
        rom[2096] = 24'b000010011011001001110001;
        rom[2097] = 24'b000001010011110010110111;
        rom[2098] = 24'b000001000011001010000100;
        rom[2099] = 24'b000001111100000100110011;
        rom[2100] = 24'b000011000000000001001010;
        rom[2101] = 24'b000010111101001010000100;
        rom[2102] = 24'b000010000011000000001011;
        rom[2103] = 24'b000001001000111000010110;
        rom[2104] = 24'b000001011100100110100111;
        rom[2105] = 24'b000010100000000100100110;
        rom[2106] = 24'b000011000101110000010000;
        rom[2107] = 24'b000010100111011001010110;
        rom[2108] = 24'b000001101000110011110111;
        rom[2109] = 24'b000001001011010100100110;
        rom[2110] = 24'b000001111011101011011011;
        rom[2111] = 24'b000010111101001010000100;
        rom[2112] = 24'b000011000010011101011010;
        rom[2113] = 24'b000010001010101110010011;
        rom[2114] = 24'b000001010001110011100100;
        rom[2115] = 24'b000001011101100011110111;
        rom[2116] = 24'b000010011000101101100001;
        rom[2117] = 24'b000011000000101000111000;
        rom[2118] = 24'b000010101001101011011000;
        rom[2119] = 24'b000001101010100101111101;
        rom[2120] = 24'b000001001010001010110110;
        rom[2121] = 24'b000001111000111010111111;
        rom[2122] = 24'b000010110010100101110111;
        rom[2123] = 24'b000010111101100110000000;
        rom[2124] = 24'b000010001011001010010000;
        rom[2125] = 24'b000001010110010010001111;
        rom[2126] = 24'b000001011100011001111000;
        rom[2127] = 24'b000010010110000100110000;
        rom[2128] = 24'b000010111101100000001001;
        rom[2129] = 24'b000010100110110110000010;
        rom[2130] = 24'b000001101010001100111000;
        rom[2131] = 24'b000001010000110011000111;
        rom[2132] = 24'b000001111000101110011110;
        rom[2133] = 24'b000010110110010100011000;
        rom[2134] = 24'b000010111010101111111011;
        rom[2135] = 24'b000010001011100110001100;
        rom[2136] = 24'b000001001110111110100101;
        rom[2137] = 24'b000001010110101110001011;
        rom[2138] = 24'b000010001110011011110100;
        rom[2139] = 24'b000010111100010110011001;
        rom[2140] = 24'b000010011110110111001000;
        rom[2141] = 24'b000001100000010001101001;
        rom[2142] = 24'b000001000100010111000000;
        rom[2143] = 24'b000001101010000010101001;
        rom[2144] = 24'b000010101000101000001000;
        rom[2145] = 24'b000010111100010110011001;
        rom[2146] = 24'b000010000111000111000100;
        rom[2147] = 24'b000001010001110101101011;
        rom[2148] = 24'b000001010011110111000101;
        rom[2149] = 24'b000010010010111010111100;
        rom[2150] = 24'b000011000100100000111011;
        rom[2151] = 24'b000010110001011011111000;
        rom[2152] = 24'b000001101100100001001110;
        rom[2153] = 24'b000001001011111010100111;
        rom[2154] = 24'b000001110011111101110111;
        rom[2155] = 24'b000010110101011111100010;
        rom[2156] = 24'b000011001110100101111001;
        rom[2157] = 24'b000010011010111101010000;
        rom[2158] = 24'b000001100011101110101000;
        rom[2159] = 24'b000001100010011111011111;
        rom[2160] = 24'b000010011110101100001111;
        rom[2161] = 24'b000011011000011100110000;
        rom[2162] = 24'b000011010010010101000111;
        rom[2163] = 24'b000010010001010101011111;
        rom[2164] = 24'b000001011101101100110110;
        rom[2165] = 24'b000010000000100100001101;
        rom[2166] = 24'b000011000110111110010111;
        rom[2167] = 24'b000011101100100101011000;
        rom[2168] = 24'b000011000111000110010001;
        rom[2169] = 24'b000010000111000100000111;
        rom[2170] = 24'b000001110001100010110100;
        rom[2171] = 24'b000010101000000001010011;
        rom[2172] = 24'b000011100100101000111010;
        rom[2173] = 24'b000011100100001110000100;
        rom[2174] = 24'b000010100111100111111011;
        rom[2175] = 24'b000001101011000011110110;
        rom[2176] = 24'b000010000001001110010111;
        rom[2177] = 24'b000010111000011111000110;
        rom[2178] = 24'b000011100101011111100000;
        rom[2179] = 24'b000011000111001000100110;
        rom[2180] = 24'b000010000110000110110111;
        rom[2181] = 24'b000001110111010001000110;
        rom[2182] = 24'b000010100101001011101011;
        rom[2183] = 24'b000011100001110001110100;
        rom[2184] = 24'b000011101001100001011010;
        rom[2185] = 24'b000010101100111001110011;
        rom[2186] = 24'b000001111000110111100100;
        rom[2187] = 24'b000010000010001011100111;
        rom[2188] = 24'b000010111111110001100001;
        rom[2189] = 24'b000011100101010000101000;
        rom[2190] = 24'b000011001011110110111000;
        rom[2191] = 24'b000010001111001101101101;
        rom[2192] = 24'b000001110001001110110110;
        rom[2193] = 24'b000010011000101010001111;
        rom[2194] = 24'b000011010111001101100111;
        rom[2195] = 24'b000011011101010101010000;
        rom[2196] = 24'b000010101101010101110000;
        rom[2197] = 24'b000001110110000001011111;
        rom[2198] = 24'b000010000001000001101000;
        rom[2199] = 24'b000010110101110100000000;
        rom[2200] = 24'b000011011101001111011001;
        rom[2201] = 24'b000011000110100101010010;
        rom[2202] = 24'b000010000111011111111000;
        rom[2203] = 24'b000001100001111000110111;
        rom[2204] = 24'b000010000100111011101110;
        rom[2205] = 24'b000011000000000101011000;
        rom[2206] = 24'b000011001011110101101011;
        rom[2207] = 24'b000010100100000000101100;
        rom[2208] = 24'b000001101100010001100101;
        rom[2209] = 24'b000001101111001000101011;
        rom[2210] = 24'b000010101001010010100100;
        rom[2211] = 24'b000011010010010100101001;
        rom[2212] = 24'b000010111100001010001000;
        rom[2213] = 24'b000001111101100100101001;
        rom[2214] = 24'b000001011010010101010000;
        rom[2215] = 24'b000010000100111001011001;
        rom[2216] = 24'b000011000001000010101000;
        rom[2217] = 24'b000011001111111000011001;
        rom[2218] = 24'b000010100110110110010100;
        rom[2219] = 24'b000001100101010111101011;
        rom[2220] = 24'b000001100111011001000101;
        rom[2221] = 24'b000010100110011100111100;
        rom[2222] = 24'b000011011000000010111011;
        rom[2223] = 24'b000011000100111101111000;
        rom[2224] = 24'b000001111101100110111110;
        rom[2225] = 24'b000001011111011100100111;
        rom[2226] = 24'b000001111101101110110111;
        rom[2227] = 24'b000010111111010000100010;
        rom[2228] = 24'b000011011010110011001001;
        rom[2229] = 24'b000010101100000011000000;
        rom[2230] = 24'b000001101011000011011000;
        rom[2231] = 24'b000001100000000011001111;
        rom[2232] = 24'b000010011110101100001111;
        rom[2233] = 24'b000011010001001000000000;
        rom[2234] = 24'b000011001011000000010111;
        rom[2235] = 24'b000010000111100100011111;
        rom[2236] = 24'b000001010110011000000110;
        rom[2237] = 24'b000001110110110011001101;
        rom[2238] = 24'b000010111000010100110111;
        rom[2239] = 24'b000011011001000011011000;
        rom[2240] = 24'b000010101110101011110001;
        rom[2241] = 24'b000001101100001101010111;
        rom[2242] = 24'b000001001111010111010100;
        rom[2243] = 24'b000010000101110101110011;
        rom[2244] = 24'b000011001100001110011010;
        rom[2245] = 24'b000011001001010111010100;
        rom[2246] = 24'b000010000111111000101011;
        rom[2247] = 24'b000001010111100001110110;
        rom[2248] = 24'b000001100001011111000111;
        rom[2249] = 24'b000010101001110101100110;
        rom[2250] = 24'b000011001111100001010000;
        rom[2251] = 24'b000010110110000010110110;
        rom[2252] = 24'b000001111001111001100111;
        rom[2253] = 24'b000001100011101111000110;
        rom[2254] = 24'b000010001100110001001011;
        rom[2255] = 24'b000011001001010111010100;
        rom[2256] = 24'b000011010001000110111010;
        rom[2257] = 24'b000010010110111011100011;
        rom[2258] = 24'b000001101010001110000100;
        rom[2259] = 24'b000001101100001101010111;
        rom[2260] = 24'b000010101001110011010001;
        rom[2261] = 24'b000011010001101110101000;
        rom[2262] = 24'b000010110101111000101000;
        rom[2263] = 24'b000001110100010110111101;
        rom[2264] = 24'b000001011000110100010110;
        rom[2265] = 24'b000010000000001111101111;
        rom[2266] = 24'b000010111001111010100111;
        rom[2267] = 24'b000011000010011110100000;
        rom[2268] = 24'b000010010100111011010000;
        rom[2269] = 24'b000001011011001010101111;
        rom[2270] = 24'b000001100001010010011000;
        rom[2271] = 24'b000010100010010010000000;
        rom[2272] = 24'b000011001100001001101001;
        rom[2273] = 24'b000010110111111011110010;
        rom[2274] = 24'b000001111011010010101000;
        rom[2275] = 24'b000001011101000000010111;
        rom[2276] = 24'b000010000010011111011110;
        rom[2277] = 24'b000011000000000101011000;
        rom[2278] = 24'b000011001011110101101011;
        rom[2279] = 24'b000010011100101011111100;
        rom[2280] = 24'b000001100111011001000101;
        rom[2281] = 24'b000001101111001000101011;
        rom[2282] = 24'b000010101001010010100100;
        rom[2283] = 24'b000011011100000101101001;
        rom[2284] = 24'b000011000011011110111000;
        rom[2285] = 24'b000010000100111001011001;
        rom[2286] = 24'b000001011111001101110000;
        rom[2287] = 24'b000001111101100100101001;
        rom[2288] = 24'b000011000011011110111000;
        rom[2289] = 24'b000011010010010100101001;
        rom[2290] = 24'b000010011101000101010100;
        rom[2291] = 24'b000001100101010111101011;
        rom[2292] = 24'b000001100010100000100101;
        rom[2293] = 24'b000010011111001000001100;
        rom[2294] = 24'b000011010000101110001011;
        rom[2295] = 24'b000010111011001100111000;
        rom[2296] = 24'b000001111011001010101110;
        rom[2297] = 24'b000001010101101011100111;
        rom[2298] = 24'b000001111101101110111000;
        rom[2299] = 24'b000010111100110100010010;
        rom[2300] = 24'b000011010011011110011001;
        rom[2301] = 24'b000010100100101110010000;
        rom[2302] = 24'b000001100001010010011000;
        rom[2303] = 24'b000001011011001010101111;
        rom[2304] = 24'b000010010100111011001111;
        rom[2305] = 24'b000011001110101011110000;
        rom[2306] = 24'b000011001000100100000111;
        rom[2307] = 24'b000010000111100100011111;
        rom[2308] = 24'b000001011011010000100110;
        rom[2309] = 24'b000001111001001111011101;
        rom[2310] = 24'b000010111111101001100111;
        rom[2311] = 24'b000011011011011111101000;
        rom[2312] = 24'b000010110011100100010001;
        rom[2313] = 24'b000001101110101001100111;
        rom[2314] = 24'b000001011110000000110100;
        rom[2315] = 24'b000010010010000011000011;
        rom[2316] = 24'b000011001001110010001010;
        rom[2317] = 24'b000011010000101100000100;
        rom[2318] = 24'b000010001111001101011011;
        rom[2319] = 24'b000001100001010010110110;
        rom[2320] = 24'b000001110000001000100111;
        rom[2321] = 24'b000010110011100110100110;
        rom[2322] = 24'b000011010100011001110000;
        rom[2323] = 24'b000010111000011111000110;
        rom[2324] = 24'b000001111100010101110111;
        rom[2325] = 24'b000001101011000011110110;
        rom[2326] = 24'b000010011011011010101011;
        rom[2327] = 24'b000011100001110001110100;
        rom[2328] = 24'b000011100111000101001010;
        rom[2329] = 24'b000010101111010110000011;
        rom[2330] = 24'b000001111000110111100100;
        rom[2331] = 24'b000010001011111100100111;
        rom[2332] = 24'b000011000111000110010001;
        rom[2333] = 24'b000011111000110010101000;
        rom[2334] = 24'b000011011111011000111000;
        rom[2335] = 24'b000010100010101111101101;
        rom[2336] = 24'b000010001110100001110110;
        rom[2337] = 24'b000010111010110101101111;
        rom[2338] = 24'b000011110110111100110111;
        rom[2339] = 24'b000011111101000100100000;
        rom[2340] = 24'b000011001010101000110000;
        rom[2341] = 24'b000010010011010100011111;
        rom[2342] = 24'b000010011001011100001000;
        rom[2343] = 24'b000011001110001110100000;
        rom[2344] = 24'b000011110101101001111001;
        rom[2345] = 24'b000011100001011100000010;
        rom[2346] = 24'b000010100100110010111000;
        rom[2347] = 24'b000010001101110101010111;
        rom[2348] = 24'b000010101011111111101110;
        rom[2349] = 24'b000011100100101101001000;
        rom[2350] = 24'b000011100100010000001011;
        rom[2351] = 24'b000010111001111110111100;
        rom[2352] = 24'b000010000010001111110101;
        rom[2353] = 24'b000010010001010100001011;
        rom[2354] = 24'b000011010000010110100100;
        rom[2355] = 24'b000011111110010001001001;
        rom[2356] = 24'b000011100011001110001000;
        rom[2357] = 24'b000010011010110111101001;
        rom[2358] = 24'b000001110010101111110000;
        rom[2359] = 24'b000010010011100010111001;
        rom[2360] = 24'b000011010010001000011000;
        rom[2361] = 24'b000011010111001101001001;
        rom[2362] = 24'b000010011101000101010100;
        rom[2363] = 24'b000001100010111011011011;
        rom[2364] = 24'b000001100000000100010101;
        rom[2365] = 24'b000010011010001111101100;
        rom[2366] = 24'b000011001011110101101011;
        rom[2367] = 24'b000010111101101001001000;
        rom[2368] = 24'b000001111101100110111110;
        rom[2369] = 24'b000001010000110011000111;
        rom[2370] = 24'b000001111000110110010111;
        rom[2371] = 24'b000010110011000011010010;
        rom[2372] = 24'b000011001100001001101001;
        rom[2373] = 24'b000010010011101000100000;
        rom[2374] = 24'b000001001011010100001000;
        rom[2375] = 24'b000001001010000100111111;
        rom[2376] = 24'b000010000011110101011111;
        rom[2377] = 24'b000011000010011110100000;
        rom[2378] = 24'b000010111100010110110111;
        rom[2379] = 24'b000001110100000010011111;
        rom[2380] = 24'b000001000000011001110110;
        rom[2381] = 24'b000001011110011000101101;
        rom[2382] = 24'b000010100100110010110111;
        rom[2383] = 24'b000011000011000101001000;
        rom[2384] = 24'b000010011011001001110001;
        rom[2385] = 24'b000001010011110010110111;
        rom[2386] = 24'b000000111011110101010100;
        rom[2387] = 24'b000001101010111111000011;
        rom[2388] = 24'b000010011101110101101010;
        rom[2389] = 24'b000010001001111000110100;
        rom[2390] = 24'b000001001111101110111011;
        rom[2391] = 24'b000000001110010010010110;
        rom[2392] = 24'b000000001001100110000111;
        rom[2393] = 24'b000001001000001011100110;
        rom[2394] = 24'b000010000011110101100000;
        rom[2395] = 24'b000010010011110111010110;
        rom[2396] = 24'b000010001010111111010111;
        rom[2397] = 24'b000010101111011010110110;
        rom[2398] = 24'b000100110010110010001011;
        rom[2399] = 24'b000111100100100100010100;
        rom[2400] = 24'b001001101000110100101010;
        rom[2401] = 24'b001010011110111100110011;
        rom[2402] = 24'b001010101010011001000100;
        rom[2403] = 24'b001011001100000111100111;
        rom[2404] = 24'b001011011101110001000001;
        rom[2405] = 24'b001010010101011000111000;
        rom[2406] = 24'b000111010011100001111000;
        rom[2407] = 24'b000100000001111101011101;
        rom[2408] = 24'b000001111111111000010110;
        rom[2409] = 24'b000001100111110101001111;
        rom[2410] = 24'b000010000001110000110111;
        rom[2411] = 24'b000001110001111010010000;
        rom[2412] = 24'b000001000001111010110000;
        rom[2413] = 24'b000000011011101100001111;
        rom[2414] = 24'b000000110101010101111000;
        rom[2415] = 24'b000001111011001110000000;
        rom[2416] = 24'b000010100111100001111001;
        rom[2417] = 24'b000010010101110000010010;
        rom[2418] = 24'b000001011011100011011000;
        rom[2419] = 24'b000001000010001001100111;
        rom[2420] = 24'b000001101010000100111110;
        rom[2421] = 24'b000010100111101010111000;
        rom[2422] = 24'b000010110011011011001011;
        rom[2423] = 24'b000001111100111100101100;
        rom[2424] = 24'b000001000101001101100101;
        rom[2425] = 24'b000001000011001100001011;
        rom[2426] = 24'b000001111111110010010100;
        rom[2427] = 24'b000010101011010000101001;
        rom[2428] = 24'b000010010010101001111000;
        rom[2429] = 24'b000001010001101000001001;
        rom[2430] = 24'b000000111000001001110000;
        rom[2431] = 24'b000001011011011001001001;
        rom[2432] = 24'b000010011100011010111000;
        rom[2433] = 24'b000010101000110100011001;
        rom[2434] = 24'b000001111000011101100100;
        rom[2435] = 24'b000000111110010011101011;
        rom[2436] = 24'b000001000010110001010101;
        rom[2437] = 24'b000001111010100000011100;
        rom[2438] = 24'b000010101110100010101011;
        rom[2439] = 24'b000010100010110010011000;
        rom[2440] = 24'b000001011000111111001110;
        rom[2441] = 24'b000000110001000011110111;
        rom[2442] = 24'b000001010110101010110111;
        rom[2443] = 24'b000010010101110000010010;
        rom[2444] = 24'b000010101110110110101001;
        rom[2445] = 24'b000001111101101010010000;
        rom[2446] = 24'b000000111111000110111000;
        rom[2447] = 24'b000000111011011011011111;
        rom[2448] = 24'b000001110101001011111111;
        rom[2449] = 24'b000010101110111100100000;
        rom[2450] = 24'b000010100011111100010111;
        rom[2451] = 24'b000001100101011000111111;
        rom[2452] = 24'b000000110100001100100110;
        rom[2453] = 24'b000001010111000011111101;
        rom[2454] = 24'b000010010011101101000111;
        rom[2455] = 24'b000010110100011011101000;
        rom[2456] = 24'b000010001010000100000001;
        rom[2457] = 24'b000001000101001001010111;
        rom[2458] = 24'b000000110110111100110100;
        rom[2459] = 24'b000001101111110111100011;
        rom[2460] = 24'b000010101010000010111010;
        rom[2461] = 24'b000010101110100000100100;
        rom[2462] = 24'b000001101101000001111011;
        rom[2463] = 24'b000000111010001110110110;
        rom[2464] = 24'b000001000001101111110111;
        rom[2465] = 24'b000010000111101010000110;
        rom[2466] = 24'b000010101010111001100000;
        rom[2467] = 24'b000010001110111110110110;
        rom[2468] = 24'b000001001101111101000111;
        rom[2469] = 24'b000000110101010110010110;
        rom[2470] = 24'b000001100101101101001011;
        rom[2471] = 24'b000010100100101111100100;
        rom[2472] = 24'b000010101010000010111010;
        rom[2473] = 24'b000001110111001100010011;
        rom[2474] = 24'b000001000011001010000100;
        rom[2475] = 24'b000001001100011110000111;
        rom[2476] = 24'b000010001100100000010001;
        rom[2477] = 24'b000010110110110111111000;
        rom[2478] = 24'b000010011111111010011000;
        rom[2479] = 24'b000001011110011000101101;
        rom[2480] = 24'b000001000000011001110110;
        rom[2481] = 24'b000001101100101101101111;
        rom[2482] = 24'b000010100110011000100111;
        rom[2483] = 24'b000010101100100000010000;
        rom[2484] = 24'b000010000001011001010000;
        rom[2485] = 24'b000001001010000100111111;
        rom[2486] = 24'b000001010010101000111000;
        rom[2487] = 24'b000010010001001100010000;
        rom[2488] = 24'b000010110001010010111001;
        rom[2489] = 24'b000010011111100001010010;
        rom[2490] = 24'b000001100000011011111000;
        rom[2491] = 24'b000000111111101101010111;
        rom[2492] = 24'b000001100000010011111110;
        rom[2493] = 24'b000010011001000001011000;
        rom[2494] = 24'b000010011101011100111011;
        rom[2495] = 24'b000001101011110110111100;
        rom[2496] = 24'b000000110110100100000101;
        rom[2497] = 24'b000000110110111110111011;
        rom[2498] = 24'b000001110001001000110100;
        rom[2499] = 24'b000010011111000011011001;
        rom[2500] = 24'b000010000001100100001000;
        rom[2501] = 24'b000000111011101001111001;
        rom[2502] = 24'b000000100010001011100000;
        rom[2503] = 24'b000000111110000110001001;
        rom[2504] = 24'b000001111010001111011000;
        rom[2505] = 24'b000010010000011001111001;
        rom[2506] = 24'b000001010110010010000100;
        rom[2507] = 24'b000000100001000000101011;
        rom[2508] = 24'b000000100101011110010101;
        rom[2509] = 24'b000001011101001101011100;
        rom[2510] = 24'b000010010011101011111011;
        rom[2511] = 24'b000001111110001010101000;
        rom[2512] = 24'b000000111110001000011110;
        rom[2513] = 24'b000000011011000101100111;
        rom[2514] = 24'b000000111110010000010111;
        rom[2515] = 24'b000010001001100011000010;
        rom[2516] = 24'b000010100010101001011001;
        rom[2517] = 24'b000001110001011101000000;
        rom[2518] = 24'b000000110101010101111000;
        rom[2519] = 24'b000000111000111111001111;
        rom[2520] = 24'b000001110101001011111111;
        rom[2521] = 24'b000010101110111100100000;
        rom[2522] = 24'b000010101101101101010111;
        rom[2523] = 24'b000001101111001001111111;
        rom[2524] = 24'b000001000111101110100110;
        rom[2525] = 24'b000001100101101101011101;
        rom[2526] = 24'b000010101100000111100111;
        rom[2527] = 24'b000011010110100111001000;
        rom[2528] = 24'b000010110001001000000001;
        rom[2529] = 24'b000001101110101001100111;
        rom[2530] = 24'b000001100010111001010100;
        rom[2531] = 24'b000010011011110100000011;
        rom[2532] = 24'b000011011010110111111010;
        rom[2533] = 24'b000011011010011101000100;
        rom[2534] = 24'b000010100111100111111011;
        rom[2535] = 24'b000001101111111100010110;
        rom[2536] = 24'b000010000110000110110111;
        rom[2537] = 24'b000011001100000001000110;
        rom[2538] = 24'b000011110001101100110000;
        rom[2539] = 24'b000011001100000001000110;
        rom[2540] = 24'b000010001010111111010111;
        rom[2541] = 24'b000001110100110100110110;
        rom[2542] = 24'b000010011011011010101011;
        rom[2543] = 24'b000011100001110001110100;
        rom[2544] = 24'b000011100010001100101010;
        rom[2545] = 24'b000010101000000001010011;
        rom[2546] = 24'b000001110001100010110100;
        rom[2547] = 24'b000001111101010011000111;
        rom[2548] = 24'b000010111101010101010001;
        rom[2549] = 24'b000011100101010000101000;
        rom[2550] = 24'b000011001110010011001000;
        rom[2551] = 24'b000010001100110001011101;
        rom[2552] = 24'b000001110001001110110110;
        rom[2553] = 24'b000010011000101010001111;
        rom[2554] = 24'b000011010100110001010111;
        rom[2555] = 24'b000011011111110001100000;
        rom[2556] = 24'b000010101000011101010000;
        rom[2557] = 24'b000001110110000001011111;
        rom[2558] = 24'b000001111100001001001000;
        rom[2559] = 24'b000010110101110100000000;
        rom[2560] = 24'b000011011111101011101001;
        rom[2561] = 24'b000011001001000001100010;
        rom[2562] = 24'b000010001110110100101000;
        rom[2563] = 24'b000001101110000110000111;
        rom[2564] = 24'b000010010110000001011110;
        rom[2565] = 24'b000011001110101110111000;
        rom[2566] = 24'b000011011100111011011011;
        rom[2567] = 24'b000010101101110001101100;
        rom[2568] = 24'b000001110011100110010101;
        rom[2569] = 24'b000001111000111001101011;
        rom[2570] = 24'b000010110101011111110100;
        rom[2571] = 24'b000011100011011010011001;
        rom[2572] = 24'b000011000011011110111000;
        rom[2573] = 24'b000010000100111001011001;
        rom[2574] = 24'b000001100001101010000000;
        rom[2575] = 24'b000010001001110001111001;
        rom[2576] = 24'b000011000101111011001000;
        rom[2577] = 24'b000011010100110000111001;
        rom[2578] = 24'b000010100100011010000100;
        rom[2579] = 24'b000001100111110011111011;
        rom[2580] = 24'b000001101001110101010101;
        rom[2581] = 24'b000010101000111001001100;
        rom[2582] = 24'b000011011100111011011011;
        rom[2583] = 24'b000011001001110110011000;
        rom[2584] = 24'b000010000100111011101110;
        rom[2585] = 24'b000001100100010101000111;
        rom[2586] = 24'b000010000101000011100111;
        rom[2587] = 24'b000011001001000001100010;
        rom[2588] = 24'b000011011111101011101001;
        rom[2589] = 24'b000010101110011111010000;
        rom[2590] = 24'b000001101101011111101000;
        rom[2591] = 24'b000001100100111011101111;
        rom[2592] = 24'b000010100001001000011111;
        rom[2593] = 24'b000011011010111001000000;
        rom[2594] = 24'b000011010100110001010111;
        rom[2595] = 24'b000010000111100100011111;
        rom[2596] = 24'b000001011101101100110110;
        rom[2597] = 24'b000001111011101011101101;
        rom[2598] = 24'b000011000010000101111000;
        rom[2599] = 24'b000011011011011111101000;
        rom[2600] = 24'b000010110001001000000001;
        rom[2601] = 24'b000001101100001101010111;
        rom[2602] = 24'b000001010100001111110100;
        rom[2603] = 24'b000010001101001010100011;
        rom[2604] = 24'b000011010011100011001010;
        rom[2605] = 24'b000011010000101100000100;
        rom[2606] = 24'b000010010001101001101011;
        rom[2607] = 24'b000001011110110110100110;
        rom[2608] = 24'b000001101101101100010111;
        rom[2609] = 24'b000010110001001010010110;
        rom[2610] = 24'b000011011011101110100000;
        rom[2611] = 24'b000010111000011111000110;
        rom[2612] = 24'b000001110101000001000111;
        rom[2613] = 24'b000001011100011010010110;
        rom[2614] = 24'b000010001100110001001011;
        rom[2615] = 24'b000011001110001111110100;
        rom[2616] = 24'b000011001110101010101010;
        rom[2617] = 24'b000010011011110100000011;
        rom[2618] = 24'b000001100101010101100100;
        rom[2619] = 24'b000001101110101001100111;
        rom[2620] = 24'b000010101110101011110001;
        rom[2621] = 24'b000011010110100111001000;
        rom[2622] = 24'b000010111111101001101000;
        rom[2623] = 24'b000001111110000111111101;
        rom[2624] = 24'b000001100010100101010110;
        rom[2625] = 24'b000010000101001000001111;
        rom[2626] = 24'b000011000001001111010111;
        rom[2627] = 24'b000011010011100100010000;
        rom[2628] = 24'b000010100110000001000000;
        rom[2629] = 24'b000001110011100101001111;
        rom[2630] = 24'b000001111110100101011000;
        rom[2631] = 24'b000011000110111001110000;
        rom[2632] = 24'b000011101110010101001001;
        rom[2633] = 24'b000011011010000111010010;
        rom[2634] = 24'b000010010110001001011000;
        rom[2635] = 24'b000001111111001011110111;
        rom[2636] = 24'b000010101011111111101110;
        rom[2637] = 24'b000011110011010110101000;
        rom[2638] = 24'b000011111010001110011011;
        rom[2639] = 24'b000011001011000100101100;
        rom[2640] = 24'b000010010011010101100101;
        rom[2641] = 24'b000010011011000101001011;
        rom[2642] = 24'b000011011010000111100100;
        rom[2643] = 24'b000100000101100101111001;
        rom[2644] = 24'b000011101100111111001000;
        rom[2645] = 24'b000010101110011001101001;
        rom[2646] = 24'b000010001011001010010000;
        rom[2647] = 24'b000010110011010010001001;
        rom[2648] = 24'b000011101111011011011000;
        rom[2649] = 24'b000011111001011000101001;
        rom[2650] = 24'b000011001001000001110100;
        rom[2651] = 24'b000010001110110111111011;
        rom[2652] = 24'b000010000111001000010101;
        rom[2653] = 24'b000011000011101111111100;
        rom[2654] = 24'b000100000011111111011011;
        rom[2655] = 24'b000011111010101011011000;
        rom[2656] = 24'b000010111010101001001110;
        rom[2657] = 24'b000010001011011001000111;
        rom[2658] = 24'b000010011101011110000111;
        rom[2659] = 24'b000011011100100011100010;
        rom[2660] = 24'b000011110000110001011001;
        rom[2661] = 24'b000010111010101100100000;
        rom[2662] = 24'b000001110100110100011000;
        rom[2663] = 24'b000001100010011111011111;
        rom[2664] = 24'b000010011100001111111111;
        rom[2665] = 24'b000011010001001000000000;
        rom[2666] = 24'b000011001000100100000111;
        rom[2667] = 24'b000010000000001111101111;
        rom[2668] = 24'b000001001111000011010110;
        rom[2669] = 24'b000001101010100101111101;
        rom[2670] = 24'b000010110101111000100111;
        rom[2671] = 24'b000011011001000011011000;
        rom[2672] = 24'b000010101100001111100001;
        rom[2673] = 24'b000001101001110001000111;
        rom[2674] = 24'b000001011001001000010100;
        rom[2675] = 24'b000010001101001010100011;
        rom[2676] = 24'b000011001001110010001010;
        rom[2677] = 24'b000011001001010111010100;
        rom[2678] = 24'b000010001010010100111011;
        rom[2679] = 24'b000001010111100001110110;
        rom[2680] = 24'b000001100011111011010111;
        rom[2681] = 24'b000010100100111101000110;
        rom[2682] = 24'b000011010001111101100000;
        rom[2683] = 24'b000010110001001010010110;
        rom[2684] = 24'b000001100110010111100111;
        rom[2685] = 24'b000001010000001101000110;
        rom[2686] = 24'b000001111011101011011011;
        rom[2687] = 24'b000010111000010001100100;
        rom[2688] = 24'b000011000000000001001010;
        rom[2689] = 24'b000010001000010010000011;
        rom[2690] = 24'b000001001100111011000100;
        rom[2691] = 24'b000001001100011110000111;
        rom[2692] = 24'b000001111000111110010001;
        rom[2693] = 24'b000010001111110011111000;
        rom[2694] = 24'b000001101010001100111000;
        rom[2695] = 24'b000000100001010110011101;
        rom[2696] = 24'b111111111001100110100110;
        rom[2697] = 24'b000000011001101101001111;
        rom[2698] = 24'b000001110011000111010111;
        rom[2699] = 24'b000010110110010001010000;
        rom[2700] = 24'b000011001010101000101111;
        rom[2701] = 24'b000011011100100011111111;
        rom[2702] = 24'b000101001011101010011000;
        rom[2703] = 24'b001000000100010010010000;
        rom[2704] = 24'b001010101000001110011001;
        rom[2705] = 24'b001011110101101010100010;
        rom[2706] = 24'b001011011011001100111000;
        rom[2707] = 24'b001010011111100111100111;
        rom[2708] = 24'b001001001101011110011110;
        rom[2709] = 24'b000111001100101000111000;
        rom[2710] = 24'b000100011100011001111011;
        rom[2711] = 24'b000001110000101111011100;
        rom[2712] = 24'b000000010001111100010101;
        rom[2713] = 24'b000000100011011100111011;
        rom[2714] = 24'b000001101110101100100100;
        rom[2715] = 24'b000010101101101100111001;
        rom[2716] = 24'b000010100011101111101000;
        rom[2717] = 24'b000001100010101101111001;
        rom[2718] = 24'b000000111111011110100000;
        rom[2719] = 24'b000001101010000010101001;
        rom[2720] = 24'b000010101101100000101000;
        rom[2721] = 24'b000010111100010110011001;
        rom[2722] = 24'b000010000010001110100100;
        rom[2723] = 24'b000001000000101111111011;
        rom[2724] = 24'b000001000111101001110101;
        rom[2725] = 24'b000010000001110101001100;
        rom[2726] = 24'b000010110101110111011011;
        rom[2727] = 24'b000010100111101010111000;
        rom[2728] = 24'b000001100000010011111110;
        rom[2729] = 24'b000000111101010001000111;
        rom[2730] = 24'b000001100000011011110111;
        rom[2731] = 24'b000010100100011001110010;
        rom[2732] = 24'b000010110110001011011001;
        rom[2733] = 24'b000010001110110000000000;
        rom[2734] = 24'b000001001011010100001000;
        rom[2735] = 24'b000001001100100001001111;
        rom[2736] = 24'b000010000110010001101111;
        rom[2737] = 24'b000011000010011110100000;
        rom[2738] = 24'b000010110010100101110111;
        rom[2739] = 24'b000001110100000010011111;
        rom[2740] = 24'b000001000111101110100110;
        rom[2741] = 24'b000001100000110100111101;
        rom[2742] = 24'b000010100100110010110111;
        rom[2743] = 24'b000011000000101000111000;
        rom[2744] = 24'b000010011000101101100001;
        rom[2745] = 24'b000001011000101011010111;
        rom[2746] = 24'b000001000101100110010100;
        rom[2747] = 24'b000010000000111101010011;
        rom[2748] = 24'b000010110011110011111010;
        rom[2749] = 24'b000010110101110101010100;
        rom[2750] = 24'b000001111011101011011011;
        rom[2751] = 24'b000001000110011100000110;
        rom[2752] = 24'b000001010111101110000111;
        rom[2753] = 24'b000010010110010011100110;
        rom[2754] = 24'b000010111110011011100000;
        rom[2755] = 24'b000010011101101000010110;
        rom[2756] = 24'b000001011111000010110111;
        rom[2757] = 24'b000001000110011100000110;
        rom[2758] = 24'b000001110001111010011011;
        rom[2759] = 24'b000010110011011001000100;
        rom[2760] = 24'b000010110001010111101010;
        rom[2761] = 24'b000001111001101000100011;
        rom[2762] = 24'b000001001000000010100100;
        rom[2763] = 24'b000001010110001111000111;
        rom[2764] = 24'b000010010011110101000001;
        rom[2765] = 24'b000010111110001100101000;
        rom[2766] = 24'b000010100010010110101000;
        rom[2767] = 24'b000001100011010001001101;
        rom[2768] = 24'b000001000101010010010110;
        rom[2769] = 24'b000001110001100110001111;
        rom[2770] = 24'b000010110010100101110111;
        rom[2771] = 24'b000010111101100110000000;
        rom[2772] = 24'b000010001000101101111111;
        rom[2773] = 24'b000001001110111101011111;
        rom[2774] = 24'b000001011001111101101000;
        rom[2775] = 24'b000010010110000100110000;
        rom[2776] = 24'b000010110110001011011001;
        rom[2777] = 24'b000010011111100001010010;
        rom[2778] = 24'b000001100010111000001000;
        rom[2779] = 24'b000001000111000010000111;
        rom[2780] = 24'b000001101110111101011110;
        rom[2781] = 24'b000010100111101010111000;
        rom[2782] = 24'b000010110011011011001011;
        rom[2783] = 24'b000010000100010001011100;
        rom[2784] = 24'b000001010001011010110101;
        rom[2785] = 24'b000001010001110101101011;
        rom[2786] = 24'b000010001011111111100100;
        rom[2787] = 24'b000010110111011101111001;
        rom[2788] = 24'b000010011001111110101000;
        rom[2789] = 24'b000001100010101101111001;
        rom[2790] = 24'b000000111111011110100000;
        rom[2791] = 24'b000001101010000010101001;
        rom[2792] = 24'b000010101000101000001000;
        rom[2793] = 24'b000010110101000001101001;
        rom[2794] = 24'b000001111111110010010100;
        rom[2795] = 24'b000001000101101000011011;
        rom[2796] = 24'b000001001010000110000101;
        rom[2797] = 24'b000010000100010001011100;
        rom[2798] = 24'b000010111010101111111011;
        rom[2799] = 24'b000010100111101010111000;
        rom[2800] = 24'b000001100010110000001110;
        rom[2801] = 24'b000000111010110100110111;
        rom[2802] = 24'b000001011011100011011000;
        rom[2803] = 24'b000010100001111101100010;
        rom[2804] = 24'b000010111011000011111001;
        rom[2805] = 24'b000010001001110111100000;
        rom[2806] = 24'b000001000110011011101000;
        rom[2807] = 24'b000001000000010011111111;
        rom[2808] = 24'b000001111010000100011111;
        rom[2809] = 24'b000010111000101101100000;
        rom[2810] = 24'b000010101011010001000111;
        rom[2811] = 24'b000001101111001001111111;
        rom[2812] = 24'b000001000010110110000110;
        rom[2813] = 24'b000001101000001001101101;
        rom[2814] = 24'b000010110001000000000111;
        rom[2815] = 24'b000011010100001010111000;
        rom[2816] = 24'b000010110001001000000001;
        rom[2817] = 24'b000001110001000101110111;
        rom[2818] = 24'b000001100010111001010100;
        rom[2819] = 24'b000010011110010000010011;
        rom[2820] = 24'b000011011111110000011010;
        rom[2821] = 24'b000011100100001110000100;
        rom[2822] = 24'b000010100010101111011011;
        rom[2823] = 24'b000001110010011000100110;
        rom[2824] = 24'b000010000011101010100111;
        rom[2825] = 24'b000011001100000001000110;
        rom[2826] = 24'b000011101111010000100000;
        rom[2827] = 24'b000011010000111001100110;
        rom[2828] = 24'b000010010010010100000111;
        rom[2829] = 24'b000001111100001001100110;
        rom[2830] = 24'b000010101100100000011011;
        rom[2831] = 24'b000011101101111111000100;
        rom[2832] = 24'b000011110000110110001010;
        rom[2833] = 24'b000010111101111111100011;
        rom[2834] = 24'b000010000101000100110100;
        rom[2835] = 24'b000010010011010001010111;
        rom[2836] = 24'b000011001011111110110001;
        rom[2837] = 24'b000011111011001110111000;
        rom[2838] = 24'b000011011010100000011000;
        rom[2839] = 24'b000010011101110111001101;
        rom[2840] = 24'b000001111111111000010110;
        rom[2841] = 24'b000010100111010011101111;
        rom[2842] = 24'b000011100000111110100111;
        rom[2843] = 24'b000011101110011011000000;
        rom[2844] = 24'b000010111011111111010000;
        rom[2845] = 24'b000010000100101010111111;
        rom[2846] = 24'b000010001010110010101000;
        rom[2847] = 24'b000011000100011101100000;
        rom[2848] = 24'b000011101011111000111001;
        rom[2849] = 24'b000011011010000111010010;
        rom[2850] = 24'b000010010110001001011000;
        rom[2851] = 24'b000001111100101111100111;
        rom[2852] = 24'b000010100111000111001110;
        rom[2853] = 24'b000011011101011000011000;
        rom[2854] = 24'b000011101001001000101011;
        rom[2855] = 24'b000010111001111110111100;
        rom[2856] = 24'b000010000010001111110101;
        rom[2857] = 24'b000010000000001110011011;
        rom[2858] = 24'b000010111111010000110100;
        rom[2859] = 24'b000011101101001011011001;
        rom[2860] = 24'b000011010010001000011000;
        rom[2861] = 24'b000010010001000110101001;
        rom[2862] = 24'b000001110010101111110000;
        rom[2863] = 24'b000010011010110111101001;
        rom[2864] = 24'b000011010111000000111000;
        rom[2865] = 24'b000011100101110110101001;
        rom[2866] = 24'b000010101011101110110100;
        rom[2867] = 24'b000001110100000001001011;
        rom[2868] = 24'b000001111010111011000101;
        rom[2869] = 24'b000010110010101010001100;
        rom[2870] = 24'b000011100001110011111011;
        rom[2871] = 24'b000011010011100111011000;
        rom[2872] = 24'b000010001001110100001110;
        rom[2873] = 24'b000001101001001101100111;
        rom[2874] = 24'b000010001100011000010111;
        rom[2875] = 24'b000011001101111010000010;
        rom[2876] = 24'b000011011111101011101001;
        rom[2877] = 24'b000010110011010111110000;
        rom[2878] = 24'b000001101011000011011000;
        rom[2879] = 24'b000001101001110100001111;
        rom[2880] = 24'b000010101010111001100000;
        rom[2881] = 24'b000011100100101010000000;
        rom[2882] = 24'b000011010100110001010111;
        rom[2883] = 24'b000010010001010101011111;
        rom[2884] = 24'b000001100101000001100110;
        rom[2885] = 24'b000001111001001111011101;
        rom[2886] = 24'b000011000100100010000111;
        rom[2887] = 24'b000011100010110100011000;
        rom[2888] = 24'b000010110110000000100001;
        rom[2889] = 24'b000001110001000101110111;
        rom[2890] = 24'b000001100000011101000100;
        rom[2891] = 24'b000010011001010111110011;
        rom[2892] = 24'b000011011000011011101010;
        rom[2893] = 24'b000011010101100100100100;
        rom[2894] = 24'b000010010110100010001011;
        rom[2895] = 24'b000001100110001011010110;
        rom[2896] = 24'b000001110111011101010111;
        rom[2897] = 24'b000010111101010111100110;
        rom[2898] = 24'b000011100000100111000000;
        rom[2899] = 24'b000011000010010000000110;
        rom[2900] = 24'b000010000001001110010111;
        rom[2901] = 24'b000001101000100111100110;
        rom[2902] = 24'b000010010110100010001011;
        rom[2903] = 24'b000011010011001000010100;
        rom[2904] = 24'b000011011111110000011010;
        rom[2905] = 24'b000010101000000001010011;
        rom[2906] = 24'b000001110001100010110100;
        rom[2907] = 24'b000001111000011010100111;
        rom[2908] = 24'b000010111000011100110001;
        rom[2909] = 24'b000011100111101100111000;
        rom[2910] = 24'b000011000110111110011000;
        rom[2911] = 24'b000010001010010101001101;
        rom[2912] = 24'b000001101110110010100110;
        rom[2913] = 24'b000010011011000110011111;
        rom[2914] = 24'b000011001101011100100111;
        rom[2915] = 24'b000011011010111001000000;
        rom[2916] = 24'b000010101010111001100000;
        rom[2917] = 24'b000001111000011101101111;
        rom[2918] = 24'b000001111100001001001000;
        rom[2919] = 24'b000010111010101100100000;
        rom[2920] = 24'b000011011101001111011001;
        rom[2921] = 24'b000011001001000001100010;
        rom[2922] = 24'b000010001100011000010111;
        rom[2923] = 24'b000001110010111110100111;
        rom[2924] = 24'b000010011010111001111110;
        rom[2925] = 24'b000011011010111100001000;
        rom[2926] = 24'b000011110000011101011011;
        rom[2927] = 24'b000011000011101111111100;
        rom[2928] = 24'b000010010101110001110101;
        rom[2929] = 24'b000010011011000101001011;
        rom[2930] = 24'b000011010111101011010100;
        rom[2931] = 24'b000100000101100101111001;
        rom[2932] = 24'b000011101111011011011000;
        rom[2933] = 24'b000010111000001010101001;
        rom[2934] = 24'b000010011110101100010000;
        rom[2935] = 24'b000010111101000011001001;
        rom[2936] = 24'b000011111110000100111000;
        rom[2937] = 24'b000100011001000111111001;
        rom[2938] = 24'b000011100110010100110100;
        rom[2939] = 24'b000010100111010010011011;
        rom[2940] = 24'b000010100001111111000101;
        rom[2941] = 24'b000011011100001010011100;
        rom[2942] = 24'b000100001101110000011011;
        rom[2943] = 24'b000011111010101011011000;
        rom[2944] = 24'b000010110101110000101110;
        rom[2945] = 24'b000010010101001010000111;
        rom[2946] = 24'b000010110101111000100111;
        rom[2947] = 24'b000011110010100001110010;
        rom[2948] = 24'b000100010000100000101001;
        rom[2949] = 24'b000011100110101001000000;
        rom[2950] = 24'b000010101100111110001000;
        rom[2951] = 24'b000010110000100111011111;
        rom[2952] = 24'b000011011011101110011111;
        rom[2953] = 24'b000100000110110101100000;
        rom[2954] = 24'b000011110110111100110111;
        rom[2955] = 24'b000010110011100000111111;
        rom[2956] = 24'b000001111101011100000110;
        rom[2957] = 24'b000010010001101001111101;
        rom[2958] = 24'b000011010000101111010111;
        rom[2959] = 24'b000011101111000001101000;
        rom[2960] = 24'b000010111111110001100001;
        rom[2961] = 24'b000001111010110110110111;
        rom[2962] = 24'b000001100010111001010100;
        rom[2963] = 24'b000010010110111011100011;
        rom[2964] = 24'b000011011000011011101010;
        rom[2965] = 24'b000011010101100100100100;
        rom[2966] = 24'b000010011000111110011011;
        rom[2967] = 24'b000001100110001011010110;
        rom[2968] = 24'b000001110101000001000111;
        rom[2969] = 24'b000010110110000010110110;
        rom[2970] = 24'b000011011011101110100000;
        rom[2971] = 24'b000010111101010111100110;
        rom[2972] = 24'b000001110111011101010111;
        rom[2973] = 24'b000001011110110110100110;
        rom[2974] = 24'b000010000111111000101011;
        rom[2975] = 24'b000011001110001111110100;
        rom[2976] = 24'b000011010011100011001010;
        rom[2977] = 24'b000010011110010000010011;
        rom[2978] = 24'b000001101010001110000100;
        rom[2979] = 24'b000001111000011010100111;
        rom[2980] = 24'b000010101110101011110001;
        rom[2981] = 24'b000011010110100111001000;
        rom[2982] = 24'b000010111101001101010111;
        rom[2983] = 24'b000001110110110011001101;
        rom[2984] = 24'b000001001010001010110110;
        rom[2985] = 24'b000001011011100111111111;
        rom[2986] = 24'b000010001011100001110111;
        rom[2987] = 24'b000010000111111000100000;
        rom[2988] = 24'b000001000110110011010000;
        rom[2989] = 24'b000000000101101101111111;
        rom[2990] = 24'b000000100100010000001000;
        rom[2991] = 24'b000010010110000100110000;
        rom[2992] = 24'b000100000110101111101001;
        rom[2993] = 24'b000101000111111110100010;
        rom[2994] = 24'b000101101111011011101000;
        rom[2995] = 24'b000111011001110111010111;
        rom[2996] = 24'b001010000000101111101110;
        rom[2997] = 24'b001100011101100011011000;
        rom[2998] = 24'b001101000100001010011011;
        rom[2999] = 24'b001011010000101001101100;
        rom[3000] = 24'b000111110111110010000101;
        rom[3001] = 24'b000100011110111010101011;
        rom[3002] = 24'b000010110011000011100100;
        rom[3003] = 24'b000010011100100111001001;
        rom[3004] = 24'b000010000001100100001000;
        rom[3005] = 24'b000001100101001010001001;
        rom[3006] = 24'b000001010111111001000000;
        rom[3007] = 24'b000010000000000000111001;
        rom[3008] = 24'b000010111100001010001000;
        rom[3009] = 24'b000011001000100011101001;
        rom[3010] = 24'b000010010101110000100100;
        rom[3011] = 24'b000001011011100110101011;
        rom[3012] = 24'b000001011101101000000101;
        rom[3013] = 24'b000010010111110011011100;
        rom[3014] = 24'b000011001001011001011011;
        rom[3015] = 24'b000010110110010100011000;
        rom[3016] = 24'b000001110001011001101110;
        rom[3017] = 24'b000001001110010110110111;
        rom[3018] = 24'b000001101111000101010111;
        rom[3019] = 24'b000010101110001010110010;
        rom[3020] = 24'b000011001100001001101001;
        rom[3021] = 24'b000010011000100001000000;
        rom[3022] = 24'b000001010010101000111000;
        rom[3023] = 24'b000001001010000100111111;
        rom[3024] = 24'b000010001000101110000000;
        rom[3025] = 24'b000011000010011110100000;
        rom[3026] = 24'b000010111001111010100111;
        rom[3027] = 24'b000001111000111010111111;
        rom[3028] = 24'b000001000010110110000110;
        rom[3029] = 24'b000001100000110100111101;
        rom[3030] = 24'b000010100111001111000111;
        rom[3031] = 24'b000011000111111101101000;
        rom[3032] = 24'b000010100000000010010001;
        rom[3033] = 24'b000001011011000111100111;
        rom[3034] = 24'b000001001111010111010100;
        rom[3035] = 24'b000010000000111101010011;
        rom[3036] = 24'b000011000010011101011010;
        rom[3037] = 24'b000011000010000010100100;
        rom[3038] = 24'b000010000011000000001011;
        rom[3039] = 24'b000001010000001101000110;
        rom[3040] = 24'b000001011100100110100111;
        rom[3041] = 24'b000010100100111101000110;
        rom[3042] = 24'b000011001010101000110000;
        rom[3043] = 24'b000010101001110101100110;
        rom[3044] = 24'b000001100110010111100111;
        rom[3045] = 24'b000001001011010100100110;
        rom[3046] = 24'b000001111011101011011011;
        rom[3047] = 24'b000010111101001010000100;
        rom[3048] = 24'b000011000100111001101010;
        rom[3049] = 24'b000010001101001010100011;
        rom[3050] = 24'b000001011011100100100100;
        rom[3051] = 24'b000001100000000000000111;
        rom[3052] = 24'b000010011011001001110001;
        rom[3053] = 24'b000011000111111101101000;
        rom[3054] = 24'b000010101001101011011000;
        rom[3055] = 24'b000001101111011110011101;
        rom[3056] = 24'b000001010011111011110110;
        rom[3057] = 24'b000010000010101011111111;
        rom[3058] = 24'b000010111110110011000111;
        rom[3059] = 24'b000011000111010111000000;
        rom[3060] = 24'b000010010010011111000000;
        rom[3061] = 24'b000001100010011111011111;
        rom[3062] = 24'b000001100110001010111000;
        rom[3063] = 24'b000010011101011001100000;
        rom[3064] = 24'b000011001100001001101001;
        rom[3065] = 24'b000010110101011111100010;
        rom[3066] = 24'b000001101111000101011000;
        rom[3067] = 24'b000001011000000111110111;
        rom[3068] = 24'b000001111101100110111110;
        rom[3069] = 24'b000010111011001100111000;
        rom[3070] = 24'b000011000010000100101011;
        rom[3071] = 24'b000010010010111010111100;
        rom[3072] = 24'b000001011011001011110101;
        rom[3073] = 24'b000001011011100110101011;
        rom[3074] = 24'b000010011101000101010100;
        rom[3075] = 24'b000011001010111111111001;
        rom[3076] = 24'b000010110100110101011000;
        rom[3077] = 24'b000001110001010111011001;
        rom[3078] = 24'b000001001110001000000000;
        rom[3079] = 24'b000001111000101100001001;
        rom[3080] = 24'b000010110111010001101000;
        rom[3081] = 24'b000011001010111111111001;
        rom[3082] = 24'b000010011000001100110100;
        rom[3083] = 24'b000001011011100110101011;
        rom[3084] = 24'b000001011000101111100101;
        rom[3085] = 24'b000010010010111010111100;
        rom[3086] = 24'b000011001001011001011011;
        rom[3087] = 24'b000010110011111000001000;
        rom[3088] = 24'b000001110001011001101110;
        rom[3089] = 24'b000001001110010110110111;
        rom[3090] = 24'b000001101100101001000111;
        rom[3091] = 24'b000010110011000011010010;
        rom[3092] = 24'b000011001100001001101001;
        rom[3093] = 24'b000010011010111101010000;
        rom[3094] = 24'b000001011100011001111000;
        rom[3095] = 24'b000001010001011001101111;
        rom[3096] = 24'b000010010010011110111111;
        rom[3097] = 24'b000011001100001111100000;
        rom[3098] = 24'b000011000011101011100111;
        rom[3099] = 24'b000010000000001111101111;
        rom[3100] = 24'b000001001111000011010110;
        rom[3101] = 24'b000001111001001111011101;
        rom[3102] = 24'b000010111101001101011000;
        rom[3103] = 24'b000011100101010000101000;
        rom[3104] = 24'b000010111101010101010001;
        rom[3105] = 24'b000001111010110110110111;
        rom[3106] = 24'b000001101111000110100100;
        rom[3107] = 24'b000010100011001000110011;
        rom[3108] = 24'b000011100010001100101010;
        rom[3109] = 24'b000011011111010101100100;
        rom[3110] = 24'b000010100010101111011011;
        rom[3111] = 24'b000001111001101101010110;
        rom[3112] = 24'b000010001101011011100111;
        rom[3113] = 24'b000011010101110010000110;
        rom[3114] = 24'b000100000000010110010000;
        rom[3115] = 24'b000011011111100011000110;
        rom[3116] = 24'b000010100000111101100111;
        rom[3117] = 24'b000010000101111010100110;
        rom[3118] = 24'b000010110001011000111011;
        rom[3119] = 24'b000011110111110000000100;
        rom[3120] = 24'b000011111111011111101010;
        rom[3121] = 24'b000011000111110000100011;
        rom[3122] = 24'b000010001001111101010100;
        rom[3123] = 24'b000010010011010001010111;
        rom[3124] = 24'b000011010000110111010001;
        rom[3125] = 24'b000011111000110010101000;
        rom[3126] = 24'b000011011100111100100111;
        rom[3127] = 24'b000010100000010011011101;
        rom[3128] = 24'b000010000111001101000110;
        rom[3129] = 24'b000010110011100000111111;
        rom[3130] = 24'b000011101010101111100111;
        rom[3131] = 24'b000011110101101111110000;
        rom[3132] = 24'b000011000000110111110000;
        rom[3133] = 24'b000010001011111111101111;
        rom[3134] = 24'b000010010110111111111000;
        rom[3135] = 24'b000011010000101010110000;
        rom[3136] = 24'b000011110101101001111001;
        rom[3137] = 24'b000011011110111111110010;
        rom[3138] = 24'b000010011101011110001000;
        rom[3139] = 24'b000010000100000100010111;
        rom[3140] = 24'b000010101110011011111110;
        rom[3141] = 24'b000011101001100101101000;
        rom[3142] = 24'b000011110000011101011011;
        rom[3143] = 24'b000011000011101111111100;
        rom[3144] = 24'b000010001110011101000101;
        rom[3145] = 24'b000010010001010100001011;
        rom[3146] = 24'b000011001011011110000100;
        rom[3147] = 24'b000011110110111100011001;
        rom[3148] = 24'b000011011011111001011000;
        rom[3149] = 24'b000010011101010011111001;
        rom[3150] = 24'b000001111100100000110000;
        rom[3151] = 24'b000010011101010011111001;
        rom[3152] = 24'b000011011011111001011000;
        rom[3153] = 24'b000011110100100000001001;
        rom[3154] = 24'b000010111100110100100100;
        rom[3155] = 24'b000010000101000110111011;
        rom[3156] = 24'b000010000100101100000101;
        rom[3157] = 24'b000010111100011011001100;
        rom[3158] = 24'b000011110010111001101011;
        rom[3159] = 24'b000011011010111100001000;
        rom[3160] = 24'b000010010110000001011110;
        rom[3161] = 24'b000001110000100010010111;
        rom[3162] = 24'b000010001110110100100111;
        rom[3163] = 24'b000011010111101011000010;
        rom[3164] = 24'b000011101110010101001001;
        rom[3165] = 24'b000010111101001000110000;
        rom[3166] = 24'b000001110111010000101000;
        rom[3167] = 24'b000001110011100101001111;
        rom[3168] = 24'b000010110010001110001111;
        rom[3169] = 24'b000011100100101010000000;
        rom[3170] = 24'b000011100000111110100111;
        rom[3171] = 24'b000010011101100010101111;
        rom[3172] = 24'b000001101100010110010110;
        rom[3173] = 24'b000010001100110001011101;
        rom[3174] = 24'b000011010101100111110111;
        rom[3175] = 24'b000011110001011101111000;
        rom[3176] = 24'b000011000111000110010001;
        rom[3177] = 24'b000010000100100111110111;
        rom[3178] = 24'b000001101111000110100100;
        rom[3179] = 24'b000010101000000001010011;
        rom[3180] = 24'b000011100010001100101010;
        rom[3181] = 24'b000011100100001110000100;
        rom[3182] = 24'b000010100111100111111011;
        rom[3183] = 24'b000001101101100000000110;
        rom[3184] = 24'b000010000011101010100111;
        rom[3185] = 24'b000011000100101100010110;
        rom[3186] = 24'b000011101100110100010000;
        rom[3187] = 24'b000011001100000001000110;
        rom[3188] = 24'b000010000011101010100111;
        rom[3189] = 24'b000001101111111100010110;
        rom[3190] = 24'b000010100000010011001011;
        rom[3191] = 24'b000011100001110001110100;
        rom[3192] = 24'b000011100111000101001010;
        rom[3193] = 24'b000010110100001110100011;
        rom[3194] = 24'b000010000010101000100100;
        rom[3195] = 24'b000010001110011000110111;
        rom[3196] = 24'b000011000111000110010001;
        rom[3197] = 24'b000011101100100101011000;
        rom[3198] = 24'b000011010011001011100111;
        rom[3199] = 24'b000010010001101001111101;
        rom[3200] = 24'b000001110011101011000110;
        rom[3201] = 24'b000010011101100010101111;
        rom[3202] = 24'b000011011100000110000111;
        rom[3203] = 24'b000011100111000110010000;
        rom[3204] = 24'b000010110111000110101111;
        rom[3205] = 24'b000001111101010110001111;
        rom[3206] = 24'b000010001000010110011000;
        rom[3207] = 24'b000010111101001000110000;
        rom[3208] = 24'b000011101011111000111001;
        rom[3209] = 24'b000011011100100011100010;
        rom[3210] = 24'b000010100111001111001000;
        rom[3211] = 24'b000010010101001010000111;
        rom[3212] = 24'b000010110101110000101110;
        rom[3213] = 24'b000011111101000111101000;
        rom[3214] = 24'b000100000110011011101011;
        rom[3215] = 24'b000011011110100110101100;
        rom[3216] = 24'b000010100100011011010101;
        rom[3217] = 24'b000010101100001010111011;
        rom[3218] = 24'b000011101011001101010100;
        rom[3219] = 24'b000100100000011100101001;
        rom[3220] = 24'b000100001111001010101000;
        rom[3221] = 24'b000011001110001000111001;
        rom[3222] = 24'b000010110010001110010000;
        rom[3223] = 24'b000011010111111001111001;
        rom[3224] = 24'b000100010110011111011000;
        rom[3225] = 24'b000100011110000000011001;
        rom[3226] = 24'b000011101000110001000100;
        rom[3227] = 24'b000010101110100111001011;
        rom[3228] = 24'b000010101011110000000101;
        rom[3229] = 24'b000011100101111011011100;
        rom[3230] = 24'b000100011001111101101011;
        rom[3231] = 24'b000100001001010100111000;
        rom[3232] = 24'b000011000100011010001110;
        rom[3233] = 24'b000010100011110011100111;
        rom[3234] = 24'b000011010000101111010111;
        rom[3235] = 24'b000100010111001001100010;
        rom[3236] = 24'b000100101000111011001001;
        rom[3237] = 24'b000011100001110000100000;
        rom[3238] = 24'b000010011011111000011000;
        rom[3239] = 24'b000010010011010100011111;
        rom[3240] = 24'b000011000011010011111111;
        rom[3241] = 24'b000011111000001100000000;
        rom[3242] = 24'b000011101010101111100111;
        rom[3243] = 24'b000010100100110111011111;
        rom[3244] = 24'b000001111000100011100110;
        rom[3245] = 24'b000010001010010101001101;
        rom[3246] = 24'b000011010000101111010111;
        rom[3247] = 24'b000011110001011101111000;
        rom[3248] = 24'b000011001011111110110001;
        rom[3249] = 24'b000010001001100000010111;
        rom[3250] = 24'b000001110011111111000100;
        rom[3251] = 24'b000010101010011101100011;
        rom[3252] = 24'b000011100100101000111010;
        rom[3253] = 24'b000011100110101010010100;
        rom[3254] = 24'b000010101010000100001011;
        rom[3255] = 24'b000001110111010001000110;
        rom[3256] = 24'b000010000110000110110111;
        rom[3257] = 24'b000011000010010000000110;
        rom[3258] = 24'b000011100111111011110000;
        rom[3259] = 24'b000011000100101100010110;
        rom[3260] = 24'b000010000011101010100111;
        rom[3261] = 24'b000001101101100000000110;
        rom[3262] = 24'b000010010110100010001011;
        rom[3263] = 24'b000011010101100100100100;
        rom[3264] = 24'b000011011101010100001010;
        rom[3265] = 24'b000010101000000001010011;
        rom[3266] = 24'b000001110001100010110100;
        rom[3267] = 24'b000001110011100010000111;
        rom[3268] = 24'b000010100111010111000001;
        rom[3269] = 24'b000011000011000101001000;
        rom[3270] = 24'b000010010110001001011000;
        rom[3271] = 24'b000001001010110110101101;
        rom[3272] = 24'b000000100111111111010110;
        rom[3273] = 24'b000000111110010100111111;
        rom[3274] = 24'b000001110011000111010111;
        rom[3275] = 24'b000010010001101001100000;
        rom[3276] = 24'b000010010010011111000000;
        rom[3277] = 24'b000010011101000101011111;
        rom[3278] = 24'b000011101100011100101000;
        rom[3279] = 24'b000110001010001101110000;
        rom[3280] = 24'b001000111010010111001001;
        rom[3281] = 24'b001010101001111110110010;
        rom[3282] = 24'b001010111001000001011000;
        rom[3283] = 24'b001010110000101101010111;
        rom[3284] = 24'b001010011001001010001110;
        rom[3285] = 24'b001001001110000010001000;
        rom[3286] = 24'b000110011101110011001011;
        rom[3287] = 24'b000011001000101000011100;
        rom[3288] = 24'b000001000000010101000101;
        rom[3289] = 24'b000000110100100010101011;
        rom[3290] = 24'b000010000111000111000100;
        rom[3291] = 24'b000011000110000111011001;
        rom[3292] = 24'b000010111100001010001000;
        rom[3293] = 24'b000010000000000000111001;
        rom[3294] = 24'b000001011100110001100000;
        rom[3295] = 24'b000010000100111001011001;
        rom[3296] = 24'b000011000011011110111000;
        rom[3297] = 24'b000011010111001101001001;
        rom[3298] = 24'b000010100001111101110100;
        rom[3299] = 24'b000001101100101100011011;
        rom[3300] = 24'b000001101100010001100101;
        rom[3301] = 24'b000010100110011100111100;
        rom[3302] = 24'b000011011100111011011011;
        rom[3303] = 24'b000011001110101110111000;
        rom[3304] = 24'b000010000100111011101110;
        rom[3305] = 24'b000001100001111000110111;
        rom[3306] = 24'b000010000010100111011000;
        rom[3307] = 24'b000011000110100101010010;
        rom[3308] = 24'b000011011101001111011001;
        rom[3309] = 24'b000010101100000011000000;
        rom[3310] = 24'b000001100110001010111000;
        rom[3311] = 24'b000001100000000011001111;
        rom[3312] = 24'b000010010100111011001111;
        rom[3313] = 24'b000011010011100100010000;
        rom[3314] = 24'b000011001101011100100111;
        rom[3315] = 24'b000010000101001000001111;
        rom[3316] = 24'b000001011011010000100110;
        rom[3317] = 24'b000001111001001111011101;
        rom[3318] = 24'b000010111000010100110111;
        rom[3319] = 24'b000011011001000011011000;
        rom[3320] = 24'b000010101110101011110001;
        rom[3321] = 24'b000001110001000101110111;
        rom[3322] = 24'b000001011110000000110100;
        rom[3323] = 24'b000010011110010000010011;
        rom[3324] = 24'b000011011000011011101010;
        rom[3325] = 24'b000011011000000000110100;
        rom[3326] = 24'b000010010110100010001011;
        rom[3327] = 24'b000001100001010010110110;
        rom[3328] = 24'b000001110101000001000111;
        rom[3329] = 24'b000010111000011111000110;
        rom[3330] = 24'b000011100000100111000000;
        rom[3331] = 24'b000010111000011111000110;
        rom[3332] = 24'b000001110010100100110111;
        rom[3333] = 24'b000001011110110110100110;
        rom[3334] = 24'b000010000111111000101011;
        rom[3335] = 24'b000011001011110011100100;
        rom[3336] = 24'b000011010001000110111010;
        rom[3337] = 24'b000010011001010111110011;
        rom[3338] = 24'b000001011011100100100100;
        rom[3339] = 24'b000001101001110001000111;
        rom[3340] = 24'b000010100111010111000001;
        rom[3341] = 24'b000011010001101110101000;
        rom[3342] = 24'b000010111000010100111000;
        rom[3343] = 24'b000001111011101011101101;
        rom[3344] = 24'b000001100010100101010110;
        rom[3345] = 24'b000010001110111001001111;
        rom[3346] = 24'b000011001111111000110111;
        rom[3347] = 24'b000011011010111001000000;
        rom[3348] = 24'b000010101000011101010000;
        rom[3349] = 24'b000001101100010000011111;
        rom[3350] = 24'b000001101111111011111000;
        rom[3351] = 24'b000010101100000011000000;
        rom[3352] = 24'b000011011000010110111001;
        rom[3353] = 24'b000010111100110100010010;
        rom[3354] = 24'b000001111011010010101000;
        rom[3355] = 24'b000001011010100100000111;
        rom[3356] = 24'b000010000111010111111110;
        rom[3357] = 24'b000011000010100001101000;
        rom[3358] = 24'b000011001110010001111011;
        rom[3359] = 24'b000010100100000000101100;
        rom[3360] = 24'b000001101001110101010101;
        rom[3361] = 24'b000001110100000001001011;
        rom[3362] = 24'b000010100110110110010100;
        rom[3363] = 24'b000011011001101001011001;
        rom[3364] = 24'b000011000001000010101000;
        rom[3365] = 24'b000010000010011101001001;
        rom[3366] = 24'b000001100100000110010000;
        rom[3367] = 24'b000010001001110001111001;
        rom[3368] = 24'b000011000011011110111000;
        rom[3369] = 24'b000011001111111000011001;
        rom[3370] = 24'b000010011000001100110100;
        rom[3371] = 24'b000001011001001010011011;
        rom[3372] = 24'b000001100100111100110101;
        rom[3373] = 24'b000010011100101011111100;
        rom[3374] = 24'b000011010011001010011011;
        rom[3375] = 24'b000010111101101001001000;
        rom[3376] = 24'b000001110110010010001110;
        rom[3377] = 24'b000001010101101011100111;
        rom[3378] = 24'b000001110011111101110111;
        rom[3379] = 24'b000010111111010000100010;
        rom[3380] = 24'b000011011010110011001001;
        rom[3381] = 24'b000010100100101110010000;
        rom[3382] = 24'b000001100110001010111000;
        rom[3383] = 24'b000001100000000011001111;
        rom[3384] = 24'b000010011110101100001111;
        rom[3385] = 24'b000011011101010101010000;
        rom[3386] = 24'b000011010100110001010111;
        rom[3387] = 24'b000010010110001101111111;
        rom[3388] = 24'b000001100111011101110110;
        rom[3389] = 24'b000010001010010101001101;
        rom[3390] = 24'b000011001110010011000111;
        rom[3391] = 24'b000011111000110010101000;
        rom[3392] = 24'b000011001110011011000001;
        rom[3393] = 24'b000010001110011000110111;
        rom[3394] = 24'b000001111011010011110100;
        rom[3395] = 24'b000010111001000111000011;
        rom[3396] = 24'b000011110101101110101010;
        rom[3397] = 24'b000011111010001100010100;
        rom[3398] = 24'b000010111101100110001011;
        rom[3399] = 24'b000010001000010110110110;
        rom[3400] = 24'b000010011110100001010111;
        rom[3401] = 24'b000011100100011011100110;
        rom[3402] = 24'b000100001010000111010000;
        rom[3403] = 24'b000011101001010100000110;
        rom[3404] = 24'b000010101000010010010111;
        rom[3405] = 24'b000010001111101011100110;
        rom[3406] = 24'b000010111011001001111011;
        rom[3407] = 24'b000011111010001100010100;
        rom[3408] = 24'b000011111111011111101010;
        rom[3409] = 24'b000011001100101001000011;
        rom[3410] = 24'b000010010011101110010100;
        rom[3411] = 24'b000010011111011110100111;
        rom[3412] = 24'b000011010101101111110001;
        rom[3413] = 24'b000011111101101011001000;
        rom[3414] = 24'b000011100100010001011000;
        rom[3415] = 24'b000010100000010011011101;
        rom[3416] = 24'b000010000100110000110110;
        rom[3417] = 24'b000010101110101000011111;
        rom[3418] = 24'b000011101000010011010111;
        rom[3419] = 24'b000011110101101111110000;
        rom[3420] = 24'b000011000000110111110000;
        rom[3421] = 24'b000010001011111111101111;
        rom[3422] = 24'b000010010100100011101000;
        rom[3423] = 24'b000011001110001110100000;
        rom[3424] = 24'b000011110101101001111001;
        rom[3425] = 24'b000011100001011100000010;
        rom[3426] = 24'b000010011101011110000111;
        rom[3427] = 24'b000010000100000100010111;
        rom[3428] = 24'b000010100100101010111110;
        rom[3429] = 24'b000011101001100101101000;
        rom[3430] = 24'b000011110010111001101011;
        rom[3431] = 24'b000011000011101111111100;
        rom[3432] = 24'b000010000111001000010101;
        rom[3433] = 24'b000010001110110111111011;
        rom[3434] = 24'b000011001001000001110100;
        rom[3435] = 24'b000011110010000011111001;
        rom[3436] = 24'b000011011001011101001000;
        rom[3437] = 24'b000010011010110111101001;
        rom[3438] = 24'b000001110111101000010000;
        rom[3439] = 24'b000010011000011011011001;
        rom[3440] = 24'b000011010100100100101000;
        rom[3441] = 24'b000011100101110110101001;
        rom[3442] = 24'b000010111010011000010100;
        rom[3443] = 24'b000001111101110010001011;
        rom[3444] = 24'b000001111111110011100101;
        rom[3445] = 24'b000010110101000110011100;
        rom[3446] = 24'b000011101001001000101011;
        rom[3447] = 24'b000011010110000011101000;
        rom[3448] = 24'b000010010011100101001110;
        rom[3449] = 24'b000001110010111110100111;
        rom[3450] = 24'b000010001100011000010111;
        rom[3451] = 24'b000011010010110010100010;
        rom[3452] = 24'b000011101011111000111001;
        rom[3453] = 24'b000010111101001000110000;
        rom[3454] = 24'b000001111001101100111000;
        rom[3455] = 24'b000001110110000001011111;
        rom[3456] = 24'b000010110010001110001111;
        rom[3457] = 24'b000011100100101010000000;
        rom[3458] = 24'b000011011110100010010111;
        rom[3459] = 24'b000010011011000110011111;
        rom[3460] = 24'b000001101100010110010110;
        rom[3461] = 24'b000010000101011100101101;
        rom[3462] = 24'b000011001001011010100111;
        rom[3463] = 24'b000011101111000001101000;
        rom[3464] = 24'b000011000111000110010001;
        rom[3465] = 24'b000010001001100000010111;
        rom[3466] = 24'b000001110011111111000100;
        rom[3467] = 24'b000010101111010110000011;
        rom[3468] = 24'b000011100100101000111010;
        rom[3469] = 24'b000011011111010101100100;
        rom[3470] = 24'b000010100111100111111011;
        rom[3471] = 24'b000001110100110100110110;
        rom[3472] = 24'b000010000011101010100111;
        rom[3473] = 24'b000011001001100100110110;
        rom[3474] = 24'b000011110001101100110000;
        rom[3475] = 24'b000011010000111001100110;
        rom[3476] = 24'b000010001101011011100111;
        rom[3477] = 24'b000001110010011000100110;
        rom[3478] = 24'b000010011101110110111011;
        rom[3479] = 24'b000011011010011101000100;
        rom[3480] = 24'b000011100111000101001010;
        rom[3481] = 24'b000010101010011101100011;
        rom[3482] = 24'b000010000000001100010100;
        rom[3483] = 24'b000010000010001011100111;
        rom[3484] = 24'b000010111101010101010001;
        rom[3485] = 24'b000011100111101100111000;
        rom[3486] = 24'b000011011000000100001000;
        rom[3487] = 24'b000010011011011010111101;
        rom[3488] = 24'b000010001100000101100110;
        rom[3489] = 24'b000010111000011001011111;
        rom[3490] = 24'b000011110100100000100111;
        rom[3491] = 24'b000011111111100000110000;
        rom[3492] = 24'b000011001101000101000000;
        rom[3493] = 24'b000010011111100001101111;
        rom[3494] = 24'b000010101100111110001000;
        rom[3495] = 24'b000011101011100001100000;
        rom[3496] = 24'b000100010000100000101001;
        rom[3497] = 24'b000011111110101111000010;
        rom[3498] = 24'b000011000100100010001000;
        rom[3499] = 24'b000010100110001111110111;
        rom[3500] = 24'b000011001011101110111110;
        rom[3501] = 24'b000100001011110001001000;
        rom[3502] = 24'b000100010000001100101011;
        rom[3503] = 24'b000011010111010001111100;
        rom[3504] = 24'b000010100001111111000101;
        rom[3505] = 24'b000010100111010010011011;
        rom[3506] = 24'b000011011111000000000100;
        rom[3507] = 24'b000100001000000010001001;
        rom[3508] = 24'b000011101100111111001000;
        rom[3509] = 24'b000010101110011001101001;
        rom[3510] = 24'b000010010010011111000000;
        rom[3511] = 24'b000011000100010111111001;
        rom[3512] = 24'b000100000101011001101000;
        rom[3513] = 24'b000100001010011110011001;
        rom[3514] = 24'b000011001001000001110100;
        rom[3515] = 24'b000010001110110111111011;
        rom[3516] = 24'b000010001100000000110101;
        rom[3517] = 24'b000010111100011011001100;
        rom[3518] = 24'b000011101001001000101011;
        rom[3519] = 24'b000011010011100111011000;
        rom[3520] = 24'b000010001100010000011110;
        rom[3521] = 24'b000001100100010101000111;
        rom[3522] = 24'b000010001001111100001000;
        rom[3523] = 24'b000011010000010110010010;
        rom[3524] = 24'b000011101011111000111001;
        rom[3525] = 24'b000010111101001000110000;
        rom[3526] = 24'b000001110111010000101000;
        rom[3527] = 24'b000001101110101100101111;
        rom[3528] = 24'b000010101000011101010000;
        rom[3529] = 24'b000011011111110001100000;
        rom[3530] = 24'b000011010010010101000111;
        rom[3531] = 24'b000010001110111001001111;
        rom[3532] = 24'b000001100000001001000110;
        rom[3533] = 24'b000001111001001111011101;
        rom[3534] = 24'b000010111010110001000111;
        rom[3535] = 24'b000011011011011111101000;
        rom[3536] = 24'b000010110001001000000001;
        rom[3537] = 24'b000001101001110001000111;
        rom[3538] = 24'b000001011110000000110100;
        rom[3539] = 24'b000010010110111011100011;
        rom[3540] = 24'b000011001110101010101010;
        rom[3541] = 24'b000011010000101100000100;
        rom[3542] = 24'b000010010100000101111011;
        rom[3543] = 24'b000001100001010010110110;
        rom[3544] = 24'b000001101101101100010111;
        rom[3545] = 24'b000010100111011001010110;
        rom[3546] = 24'b000010111110011011100000;
        rom[3547] = 24'b000010010001011011000110;
        rom[3548] = 24'b000001001001000100100111;
        rom[3549] = 24'b000000100110101100110110;
        rom[3550] = 24'b000000111110101001001011;
        rom[3551] = 24'b000001110001011110010100;
        rom[3552] = 24'b000010001100101111111010;
        rom[3553] = 24'b000010000011011001100011;
        rom[3554] = 24'b000010001110110101110100;
        rom[3555] = 24'b000011100011110101100111;
        rom[3556] = 24'b000110000101100001110001;
        rom[3557] = 24'b001000110011101110111000;
        rom[3558] = 24'b001010010001111101011000;
        rom[3559] = 24'b001010100000111111111101;
        rom[3560] = 24'b001010100010110000010110;
        rom[3561] = 24'b001010010110111010011111;
        rom[3562] = 24'b001000111110000110010111;
        rom[3563] = 24'b000110001101000111010000;
        rom[3564] = 24'b000011001010101000110000;
        rom[3565] = 24'b000001000101001100011111;
        rom[3566] = 24'b000000110010111001101000;
        rom[3567] = 24'b000001110011111001010000;
        rom[3568] = 24'b000010101110110110101001;
        rom[3569] = 24'b000010101001010010010010;
        rom[3570] = 24'b000001110001100001101000;
        rom[3571] = 24'b000001010101101011100111;
        rom[3572] = 24'b000001111011001010101110;
        rom[3573] = 24'b000010111011001100111000;
        rom[3574] = 24'b000011000010000100101011;
        rom[3575] = 24'b000010001001001001111100;
        rom[3576] = 24'b000001011000101111100101;
        rom[3577] = 24'b000001011001001010011011;
        rom[3578] = 24'b000010010101110000100100;
        rom[3579] = 24'b000011000110000111011001;
        rom[3580] = 24'b000010110010011001001000;
        rom[3581] = 24'b000001111000101100001001;
        rom[3582] = 24'b000001010101011100110000;
        rom[3583] = 24'b000001111101100100101001;
        rom[3584] = 24'b000010110100110101011000;
        rom[3585] = 24'b000011001000100011101001;
        rom[3586] = 24'b000010010101110000100100;
        rom[3587] = 24'b000001100000011111001011;
        rom[3588] = 24'b000001011101101000000101;
        rom[3589] = 24'b000010011010001111101100;
        rom[3590] = 24'b000011001001011001011011;
        rom[3591] = 24'b000010110110010100011000;
        rom[3592] = 24'b000001110011110101111110;
        rom[3593] = 24'b000001001011111010100111;
        rom[3594] = 24'b000001101100101001000111;
        rom[3595] = 24'b000010101110001010110010;
        rom[3596] = 24'b000011000010011000101001;
        rom[3597] = 24'b000010011000100001000000;
        rom[3598] = 24'b000001010101000101001000;
        rom[3599] = 24'b000001001010000100111111;

        end
        
        always @(posedge(clk))
            begin
                if(reset)
                    begin
                        data_out <= 24'b0;
                        i <= 16'b0;
                        counter <= 20'b0;
                    end
                else
                    begin
                        if(counter == 20'd360000)
                            begin
                                data_out <= rom[i];
                                counter <= 20'b0;
                                if(i == 3599) i <= 0;
                                else i <= i + 1;
                            end
                        else counter <= counter + 20'd1;
                    end
            end
            
endmodule
